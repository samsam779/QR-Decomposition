`resetall
`timescale 1ns/1ps
module QR_Engine (
    i_clk,
    i_rst,
    i_trig,
    i_data,
    o_rd_vld,
    o_last_data,
    o_y_hat,
    o_r
);

// IO description
input          i_clk;
input          i_rst;
input          i_trig;
input  [ 47:0] i_data;
output         o_rd_vld;
output         o_last_data;
output [159:0] o_y_hat;
output [319:0] o_r;

//input related
reg [4:0] cnt_r,cnt_w;
reg signed [11:0] real_h_r [0:3][0:3];
reg signed [11:0] real_h_w [0:3][0:3];
reg signed [11:0] imag_h_r [0:3][0:3];
reg signed [11:0] imag_h_w [0:3][0:3];

// reg signed [11:0] real_h_hold_r [0:3][0:3];
// reg signed [11:0] real_h_hold_w [0:3][0:3];
// reg signed [11:0] imag_h_hold_r [0:3][0:3];
// reg signed [11:0] imag_h_hold_w [0:3][0:3];
reg signed [11:0] real_h_hold1_r, real_h_hold1_w;
reg signed [11:0] real_h_hold2_r [0:1];
reg signed [11:0] real_h_hold2_w [0:1];
reg signed [11:0] real_h_hold3_r [0:3];
reg signed [11:0] real_h_hold3_w [0:3];
reg signed [11:0] imag_h_hold1_r, imag_h_hold1_w;
reg signed [11:0] imag_h_hold2_r [0:1];
reg signed [11:0] imag_h_hold2_w [0:1];
reg signed [11:0] imag_h_hold3_r [0:3];
reg signed [11:0] imag_h_hold3_w [0:3];

reg signed [9:0] real_origin_y_r [0:3];
reg signed [9:0] real_origin_y_w [0:3];
reg signed [9:0] imag_origin_y_r [0:3];
reg signed [9:0] imag_origin_y_w [0:3];

reg signed [9:0] imag_origin_y_hold_w [0:3];
reg signed [9:0] imag_origin_y_hold_r [0:3];
reg signed [9:0] real_origin_y_hold_w [0:3];
reg signed [9:0] real_origin_y_hold_r [0:3];

//output related
reg [319:0] o_r_r, o_r_w; //{r44, r34, r24, r14, r33, r23, r13, r22, r12, r11}
reg [159:0] o_y_hat_r, o_y_hat_w;
reg o_rd_vld_r, o_rd_vld_w;
reg o_last_data_r, o_last_data_w;

reg [1:0] count_2_w,count_2_r;
reg [3:0] cnt_out_r,cnt_out_w;

reg [99:0] o_r_hold_w,o_r_hold_r;

//integer 
integer i, j;


//continuous assignment
assign o_r = o_r_r;
assign o_y_hat = o_y_hat_r;
assign o_rd_vld = o_rd_vld_r;
assign o_last_data = o_last_data_r;

wire signed [22:0] mul8_result [0:7];//{2,44}
reg [21:0] square_w [0:7];
reg [11:0] square_r [0:7];
wire [23:0] vec,vec2,vec3,vec4;
wire signed [11:0] mul8 [0:1][0:7];

assign vec = (cnt_r == 5'd16)?{imag_h_r[0][0],real_h_r[0][0]} :(cnt_r == 5'd3)?{imag_h_r[0][1],real_h_r[0][1]} :(cnt_r == 5'd10)?{imag_h_r[0][2],real_h_r[0][2]}:(cnt_r == 5'd17)?{imag_h_r[0][3],real_h_r[0][3]}:0;
assign vec2 = (cnt_r == 5'd16)?{imag_h_r[1][0],real_h_r[1][0]} :(cnt_r == 5'd3)?{imag_h_r[1][1],real_h_r[1][1]}:(cnt_r == 5'd10)?{imag_h_r[1][2],real_h_r[1][2]} :(cnt_r == 5'd17)?{imag_h_r[1][3],real_h_r[1][3]}:0;
assign vec3 = (cnt_r == 5'd16)?{imag_h_r[2][0],real_h_r[2][0]} :(cnt_r == 5'd3)?{imag_h_r[2][1],real_h_r[2][1]} :(cnt_r == 5'd10)?{imag_h_r[2][2],real_h_r[2][2]} :(cnt_r == 5'd17)?{imag_h_r[2][3],real_h_r[2][3]}:0;
assign vec4 = (cnt_r == 5'd16)?{imag_h_r[3][0],real_h_r[3][0]} :(cnt_r == 5'd3)?{imag_h_r[3][1],real_h_r[3][1]} :(cnt_r == 5'd10)?{imag_h_r[3][2],real_h_r[3][2]} :(cnt_r == 5'd17)?{imag_h_r[3][3],real_h_r[3][3]}:0;

reg [14:0] mul_add;//{5,44}
wire [21:0] sqrt_val;//{3,19}
wire [21:0] div_val_wire;//{4,18}
reg [21:0] div_val_w;
reg [21:0] div_val_r;
// assign square_wire[0] = $signed(vec[23:12])*$signed(vec[23:12]);// {S1.22}*{S1.22} = {2.44}
// assign square_wire[1] = $signed(vec[11:0])*$signed(vec[11:0]);// {s1,10}*{s1,10} = {2,20}
// assign square_wire[2] = $signed(vec2[23:12])*$signed(vec2[23:12]);
// assign square_wire[3] = $signed(vec2[11:0])*$signed(vec2[11:0]);
// assign square_wire[4] = $signed(vec3[23:12])*$signed(vec3[23:12]);
// assign square_wire[5] = $signed(vec3[11:0])*$signed(vec3[11:0]);
// assign square_wire[6] = $signed(vec4[23:12])*$signed(vec4[23:12]);
// assign square_wire[7] = $signed(vec4[11:0])*$signed(vec4[11:0]);

// assign mul_add = ((square_r[0] + square_r[1]) + (square_r[2] + square_r[3])) + ((square_r[4] + square_r[5]) + (square_r[6] + square_r[7]));
square_root_relate s1(.sum(mul_add),.sqrt_val(sqrt_val),.div_val(div_val_wire));

reg [39:0] q_r [0:3];
// reg [39:0] q4_r [0:3];
reg [39:0] q_w [0:3];
reg [39:0] q4_w [0:3];



wire [47:0] mul_in1 [0:3];
wire [39:0] mul_output_wire [0:3];
reg [39:0] mul_output_w [0:3];
reg [39:0] mul_output_r [0:3];
wire [39:0] mul_output_add;
wire signed [19:0] mul_imag,mul_real;
assign mul_in1[0] = (cnt_r == 5'd19)?{imag_h_r[0][1],12'd0,real_h_r[0][1],12'd0}:(cnt_r == 5'd0||cnt_r == 5'd6)?{imag_h_r[0][2],12'd0,real_h_r[0][2],12'd0}:(cnt_r == 5'd1)?{imag_h_w[0][3],12'd0,real_h_w[0][3],12'd0}:(cnt_r == 5'd7||cnt_r == 5'd13)?{imag_h_r[0][3],12'd0,real_h_r[0][3],12'd0}:0;
assign mul_in1[1] = (cnt_r == 5'd19)?{imag_h_r[1][1],12'd0,real_h_r[1][1],12'd0}:(cnt_r == 5'd0||cnt_r == 5'd6)?{imag_h_r[1][2],12'd0,real_h_r[1][2],12'd0}:(cnt_r == 5'd1)?{imag_h_w[1][3],12'd0,real_h_w[1][3],12'd0}:(cnt_r == 5'd7||cnt_r == 5'd13)?{imag_h_r[1][3],12'd0,real_h_r[1][3],12'd0}:0;
assign mul_in1[2] = (cnt_r == 5'd19)?{imag_h_r[2][1],12'd0,real_h_r[2][1],12'd0}:(cnt_r == 5'd0||cnt_r == 5'd6)?{imag_h_r[2][2],12'd0,real_h_r[2][2],12'd0}:(cnt_r == 5'd1)?{imag_h_w[2][3],12'd0,real_h_w[2][3],12'd0}:(cnt_r == 5'd7||cnt_r == 5'd13)?{imag_h_r[2][3],12'd0,real_h_r[2][3],12'd0}:0;
assign mul_in1[3] = (cnt_r == 5'd19)?{imag_h_r[3][1],12'd0,real_h_r[3][1],12'd0}:(cnt_r == 5'd0||cnt_r == 5'd6)?{imag_h_r[3][2],12'd0,real_h_r[3][2],12'd0}:(cnt_r == 5'd1)?{imag_h_w[3][3],12'd0,real_h_w[3][3],12'd0}:(cnt_r == 5'd7||cnt_r == 5'd13)?{imag_h_r[3][3],12'd0,real_h_r[3][3],12'd0}:0;
complex_mul_48_40 m1(.complex_in1(mul_in1[0]),.complex_in2({(~q_r[0][39:20])+20'd1,q_r[0][19:0]}),.output_data(mul_output_wire[0]));
complex_mul_48_40 m2(.complex_in1(mul_in1[1]),.complex_in2({(~q_r[1][39:20])+20'd1,q_r[1][19:0]}),.output_data(mul_output_wire[1]));
complex_mul_48_40 m3(.complex_in1(mul_in1[2]),.complex_in2({(~q_r[2][39:20])+20'd1,q_r[2][19:0]}),.output_data(mul_output_wire[2]));
complex_mul_48_40 m4(.complex_in1(mul_in1[3]),.complex_in2({(~q_r[3][39:20])+20'd1,q_r[3][19:0]}),.output_data(mul_output_wire[3]));
assign mul_imag = ($signed(mul_output_r[0][39:20]) + $signed(mul_output_r[1][39:20])) + ($signed(mul_output_r[2][39:20])+ $signed(mul_output_r[3][39:20]));
assign mul_real = ($signed(mul_output_r[0][19:0]) + $signed(mul_output_r[1][19:0])) + ($signed(mul_output_r[2][19:0])+ $signed(mul_output_r[3][19:0]));
// assign mul_output_add = {($signed(mul_output_r[0][39:20]) + $signed(mul_output_r[1][39:20])) + ($signed(mul_output_r[2][39:20])+ $signed(mul_output_r[3][39:20])),($signed(mul_output_r[0][19:0]) + $signed(mul_output_r[1][19:0])) + ($signed(mul_output_r[2][19:0])+ $signed(mul_output_r[3][19:0]))}; 
assign mul_output_add = {mul_imag,mul_real};
wire [39:0] mul_in2;
// wire [47:0] mul_output2_wire [0:3];
reg [23:0] mul_output2_w [0:3];
reg [23:0] mul_output2_r [0:3];
assign mul_in2 = (cnt_r == 5'd1)?o_r_hold_r[59:20]:(cnt_r == 5'd2)?o_r_hold_r[99:60]:(cnt_r == 5'd3)?o_r_r[219:180]:(cnt_r == 5'd8)?o_r_r[159:120]:(cnt_r == 5'd9)?o_r_r[259:220]:(cnt_r == 5'd15)?o_r_r[299:260]:0;

// complex_mul_40_40 m5(.complex_in1(mul_in2),.complex_in2({(q_r[0][39:20]),q_r[0][19:0]}),.output_data(mul_output2_wire[0]));
// complex_mul_40_40 m6(.complex_in1(mul_in2),.complex_in2({(q_r[1][39:20]),q_r[1][19:0]}),.output_data(mul_output2_wire[1]));
// complex_mul_40_40 m7(.complex_in1(mul_in2),.complex_in2({(q_r[2][39:20]),q_r[2][19:0]}),.output_data(mul_output2_wire[2]));
// complex_mul_40_40 m8(.complex_in1(mul_in2),.complex_in2({(q_r[3][39:20]),q_r[3][19:0]}),.output_data(mul_output2_wire[3]));

// wire [39:0] q_output_wire[0:3];
reg [39:0] q_output_w [0:3];
reg [39:0] q_output_r[0:3];
wire [39:0] q_in [0:3];
assign q_in[0] = (cnt_r == 5'd0)? {~q_output_r[0][39:20]+20'd1,q_output_r[0][19:0]}:{~q_r[0][39:20]+20'd1,q_r[0][19:0]};
assign q_in[1] = (cnt_r == 5'd0)? {~q_output_r[1][39:20]+20'd1,q_output_r[1][19:0]}:{~q_r[1][39:20]+20'd1,q_r[1][19:0]};
assign q_in[2] = (cnt_r == 5'd0)? {~q_output_r[2][39:20]+20'd1,q_output_r[2][19:0]}:{~q_r[2][39:20]+20'd1,q_r[2][19:0]};
assign q_in[3] = (cnt_r == 5'd0)? {~q_output_r[3][39:20]+20'd1,q_output_r[3][19:0]}:{~q_r[3][39:20]+20'd1,q_r[3][19:0]};
//final y hat calculate
wire [19:0] y_h_real,y_h_imag;

wire [39:0] y_and_mul2_in1 [0:3];
wire [39:0] y_and_mul2_in2 [0:3];
wire [31:0] y_and_mul2_out_wire [0:3];
assign y_and_mul2_in1[0] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?mul_in2:({{2{imag_origin_y_r[0][9]}},imag_origin_y_r[0],8'd0,{2{real_origin_y_r[0][9]}},real_origin_y_r[0],8'd0});
assign y_and_mul2_in1[1] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?mul_in2:({{2{imag_origin_y_r[1][9]}},imag_origin_y_r[1],8'd0,{2{real_origin_y_r[1][9]}},real_origin_y_r[1],8'd0});
assign y_and_mul2_in1[2] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?mul_in2:({{2{imag_origin_y_r[2][9]}},imag_origin_y_r[2],8'd0,{2{real_origin_y_r[2][9]}},real_origin_y_r[2],8'd0});
assign y_and_mul2_in1[3] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?mul_in2:({{2{imag_origin_y_r[3][9]}},imag_origin_y_r[3],8'd0,{2{real_origin_y_r[3][9]}},real_origin_y_r[3],8'd0});
assign y_and_mul2_in2[0] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?{(q_r[0][39:20]),q_r[0][19:0]}:q_in[0];
assign y_and_mul2_in2[1] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?{(q_r[1][39:20]),q_r[1][19:0]}:q_in[1];
assign y_and_mul2_in2[2] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?{(q_r[2][39:20]),q_r[2][19:0]}:q_in[2];
assign y_and_mul2_in2[3] = (cnt_r == 5'd1||cnt_r == 5'd2||cnt_r == 5'd3||cnt_r == 5'd8||cnt_r == 5'd9||cnt_r == 5'd15)?{(q_r[3][39:20]),q_r[3][19:0]}:q_in[3];
complex_mul_40_40 m5(.complex_in1(y_and_mul2_in1[0]),.complex_in2(y_and_mul2_in2[0]),.output_data(y_and_mul2_out_wire[0]));
complex_mul_40_40 m6(.complex_in1(y_and_mul2_in1[1]),.complex_in2(y_and_mul2_in2[1]),.output_data(y_and_mul2_out_wire[1]));
complex_mul_40_40 m7(.complex_in1(y_and_mul2_in1[2]),.complex_in2(y_and_mul2_in2[2]),.output_data(y_and_mul2_out_wire[2]));
complex_mul_40_40 m8(.complex_in1(y_and_mul2_in1[3]),.complex_in2(y_and_mul2_in2[3]),.output_data(y_and_mul2_out_wire[3]));
// complex_mul_48_40 m24(.complex_in1({imag_origin_y_r[0],14'd0,real_origin_y_r[0],14'd0}),.complex_in2(q_in[0]),.output_data(q_output_wire[0]));
// complex_mul_48_40 m25(.complex_in1({imag_origin_y_r[1],14'd0,real_origin_y_r[1],14'd0}),.complex_in2(q_in[1]),.output_data(q_output_wire[1]));
// complex_mul_48_40 m26(.complex_in1({imag_origin_y_r[2],14'd0,real_origin_y_r[2],14'd0}),.complex_in2(q_in[2]),.output_data(q_output_wire[2]));
// complex_mul_48_40 m27(.complex_in1({imag_origin_y_r[3],14'd0,real_origin_y_r[3],14'd0}),.complex_in2(q_in[3]),.output_data(q_output_wire[3]));
assign y_h_real = ($signed(q_output_r[0][19:0])+$signed(q_output_r[1][19:0]))+($signed(q_output_r[2][19:0])+$signed(q_output_r[3][19:0]));
assign y_h_imag = ($signed(q_output_r[0][39:20])+$signed(q_output_r[1][39:20]))+($signed(q_output_r[2][39:20])+$signed(q_output_r[3][39:20]));
wire signed [11:0] h_cal [0:7];
wire signed [11:0] h_result [0:7];
assign h_cal[0] = (cnt_r == 5'd16)?real_h_r[0][3]:(cnt_r == 5'd2)?real_h_r[0][1]:(cnt_r == 5'd3)?real_h_r[0][2]:(cnt_r == 5'd4)?real_h_r[0][3]:(cnt_r == 5'd9)?real_h_r[0][2]:(cnt_r == 5'd10)?real_h_r[0][3]:0;
assign h_cal[1] = (cnt_r == 5'd16)?real_h_r[1][3]:(cnt_r == 5'd2)?real_h_r[1][1]:(cnt_r == 5'd3)?real_h_r[1][2]:(cnt_r == 5'd4)?real_h_r[1][3]:(cnt_r == 5'd9)?real_h_r[1][2]:(cnt_r == 5'd10)?real_h_r[1][3]:0;
assign h_cal[2] = (cnt_r == 5'd16)?real_h_r[2][3]:(cnt_r == 5'd2)?real_h_r[2][1]:(cnt_r == 5'd3)?real_h_r[2][2]:(cnt_r == 5'd4)?real_h_r[2][3]:(cnt_r == 5'd9)?real_h_r[2][2]:(cnt_r == 5'd10)?real_h_r[2][3]:0;
assign h_cal[3] = (cnt_r == 5'd16)?real_h_r[3][3]:(cnt_r == 5'd2)?real_h_r[3][1]:(cnt_r == 5'd3)?real_h_r[3][2]:(cnt_r == 5'd4)?real_h_r[3][3]:(cnt_r == 5'd9)?real_h_r[3][2]:(cnt_r == 5'd10)?real_h_r[3][3]:0;
assign h_cal[4] = (cnt_r == 5'd16)?imag_h_r[0][3]:(cnt_r == 5'd2)?imag_h_r[0][1]:(cnt_r == 5'd3)?imag_h_r[0][2]:(cnt_r == 5'd4)?imag_h_r[0][3]:(cnt_r == 5'd9)?imag_h_r[0][2]:(cnt_r == 5'd10)?imag_h_r[0][3]:0;
assign h_cal[5] = (cnt_r == 5'd16)?imag_h_r[1][3]:(cnt_r == 5'd2)?imag_h_r[1][1]:(cnt_r == 5'd3)?imag_h_r[1][2]:(cnt_r == 5'd4)?imag_h_r[1][3]:(cnt_r == 5'd9)?imag_h_r[1][2]:(cnt_r == 5'd10)?imag_h_r[1][3]:0;
assign h_cal[6] = (cnt_r == 5'd16)?imag_h_r[2][3]:(cnt_r == 5'd2)?imag_h_r[2][1]:(cnt_r == 5'd3)?imag_h_r[2][2]:(cnt_r == 5'd4)?imag_h_r[2][3]:(cnt_r == 5'd9)?imag_h_r[2][2]:(cnt_r == 5'd10)?imag_h_r[2][3]:0;
assign h_cal[7] = (cnt_r == 5'd16)?imag_h_r[3][3]:(cnt_r == 5'd2)?imag_h_r[3][1]:(cnt_r == 5'd3)?imag_h_r[3][2]:(cnt_r == 5'd4)?imag_h_r[3][3]:(cnt_r == 5'd9)?imag_h_r[3][2]:(cnt_r == 5'd10)?imag_h_r[3][3]:0;
assign h_result[0] = h_cal[0] - $signed(mul_output2_r[0][11:0]);//h3(1)
assign h_result[1] = h_cal[1] - $signed(mul_output2_r[1][11:0]);
assign h_result[2] = h_cal[2] - $signed(mul_output2_r[2][11:0]);
assign h_result[3] = h_cal[3] - $signed(mul_output2_r[3][11:0]);
assign h_result[4] = h_cal[4] - $signed(mul_output2_r[0][23:12]);
assign h_result[5] = h_cal[5] - $signed(mul_output2_r[1][23:12]);
assign h_result[6] = h_cal[6] - $signed(mul_output2_r[2][23:12]);
assign h_result[7] = h_cal[7] - $signed(mul_output2_r[3][23:12]);

// wire signed [33:0] q_imag_tmp[0:3];//{s5,40}
// wire signed [33:0] q_real_tmp[0:3];//{s5,40}
wire signed [11:0] h_for_q_tmp[0:7];
assign h_for_q_tmp[0] = (cnt_r==5'd18)?imag_h_r[0][0]:(cnt_r==5'd19)?imag_h_r[0][3]:(cnt_r==5'd5)?imag_h_r[0][1]:(cnt_r==5'd12)?imag_h_r[0][2]:0;
assign h_for_q_tmp[1] = (cnt_r==5'd18)?imag_h_r[1][0]:(cnt_r==5'd19)?imag_h_r[1][3]:(cnt_r==5'd5)?imag_h_r[1][1]:(cnt_r==5'd12)?imag_h_r[1][2]:0;
assign h_for_q_tmp[2] = (cnt_r==5'd18)?imag_h_r[2][0]:(cnt_r==5'd19)?imag_h_r[2][3]:(cnt_r==5'd5)?imag_h_r[2][1]:(cnt_r==5'd12)?imag_h_r[2][2]:0;
assign h_for_q_tmp[3] = (cnt_r==5'd18)?imag_h_r[3][0]:(cnt_r==5'd19)?imag_h_r[3][3]:(cnt_r==5'd5)?imag_h_r[3][1]:(cnt_r==5'd12)?imag_h_r[3][2]:0;
assign h_for_q_tmp[4] = (cnt_r==5'd18)?real_h_r[0][0]:(cnt_r==5'd19)?real_h_r[0][3]:(cnt_r==5'd5)?real_h_r[0][1]:(cnt_r==5'd12)?real_h_r[0][2]:0;
assign h_for_q_tmp[5] = (cnt_r==5'd18)?real_h_r[1][0]:(cnt_r==5'd19)?real_h_r[1][3]:(cnt_r==5'd5)?real_h_r[1][1]:(cnt_r==5'd12)?real_h_r[1][2]:0;
assign h_for_q_tmp[6] = (cnt_r==5'd18)?real_h_r[2][0]:(cnt_r==5'd19)?real_h_r[2][3]:(cnt_r==5'd5)?real_h_r[2][1]:(cnt_r==5'd12)?real_h_r[2][2]:0;
assign h_for_q_tmp[7] = (cnt_r==5'd18)?real_h_r[3][0]:(cnt_r==5'd19)?real_h_r[3][3]:(cnt_r==5'd5)?real_h_r[3][1]:(cnt_r==5'd12)?real_h_r[3][2]:0;
// assign q_imag_tmp[0] = $signed({1'b0,div_val_r}) * h_for_q_tmp[0]; //{s4,18}*{s1,10}
// assign q_imag_tmp[1] = $signed({1'b0,div_val_r}) * h_for_q_tmp[1];
// assign q_imag_tmp[2] = $signed({1'b0,div_val_r}) * h_for_q_tmp[2];
// assign q_imag_tmp[3] = $signed({1'b0,div_val_r}) * h_for_q_tmp[3];
// assign q_real_tmp[0] = $signed({1'b0,div_val_r}) * h_for_q_tmp[4];
// assign q_real_tmp[1] = $signed({1'b0,div_val_r}) * h_for_q_tmp[5];
// assign q_real_tmp[2] = $signed({1'b0,div_val_r}) * h_for_q_tmp[6];
// assign q_real_tmp[3] = $signed({1'b0,div_val_r}) * h_for_q_tmp[7];
assign mul8[0][0] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec[23:12]:{1'b0,div_val_r[21:11]};
assign mul8[0][1] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec[11:0]:{1'b0,div_val_r[21:11]};
assign mul8[0][2] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec2[23:12]:{1'b0,div_val_r[21:11]};
assign mul8[0][3] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec2[11:0]:{1'b0,div_val_r[21:11]};
assign mul8[0][4] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec3[23:12]:{1'b0,div_val_r[21:11]}; 
assign mul8[0][5] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec3[11:0]:{1'b0,div_val_r[21:11]};
assign mul8[0][6] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec4[23:12]:{1'b0,div_val_r[21:11]};
assign mul8[0][7] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec4[11:0]:{1'b0,div_val_r[21:11]};
assign mul8[1][0] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec[23:12]:h_for_q_tmp[0];
assign mul8[1][1] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec[11:0]:h_for_q_tmp[1];
assign mul8[1][2] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec2[23:12]:h_for_q_tmp[2];
assign mul8[1][3] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec2[11:0]:h_for_q_tmp[3];
assign mul8[1][4] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec3[23:12]:h_for_q_tmp[4]; 
assign mul8[1][5] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec3[11:0]:h_for_q_tmp[5]; 
assign mul8[1][6] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec4[23:12]:h_for_q_tmp[6];
assign mul8[1][7] = (cnt_r==5'd16||cnt_r==5'd3||cnt_r==5'd10||cnt_r==5'd17)?vec4[11:0]:h_for_q_tmp[7];
assign mul8_result[0] = mul8[0][0]*mul8[1][0]; //{s1,10}*{s1,10}={}
assign mul8_result[1] = mul8[0][1]*mul8[1][1];
assign mul8_result[2] = mul8[0][2]*mul8[1][2];
assign mul8_result[3] = mul8[0][3]*mul8[1][3];
assign mul8_result[4] = mul8[0][4]*mul8[1][4];
assign mul8_result[5] = mul8[0][5]*mul8[1][5];
assign mul8_result[6] = mul8[0][6]*mul8[1][6];
assign mul8_result[7] = mul8[0][7]*mul8[1][7];

always @(*) begin
    //default
    for(i=0;i<4;i=i+1)begin
        for(j=0;j<4;j=j+1)begin
            real_h_w[i][j] = real_h_r[i][j];
            imag_h_w[i][j] = imag_h_r[i][j];
            // real_h_hold_w[i][j] = real_h_hold_r[i][j];
            // imag_h_hold_w[i][j] = imag_h_hold_r[i][j];
        end
        real_origin_y_w[i] = real_origin_y_r[i];
        imag_origin_y_w[i] = imag_origin_y_r[i];
        q_w[i] = q_r[i];
        q4_w[i] = 0;

        imag_origin_y_hold_w[i] = imag_origin_y_hold_r[i];
        real_origin_y_hold_w[i] = real_origin_y_hold_r[i];
        real_h_hold3_w[i] = real_h_hold3_r[i];
        imag_h_hold3_w[i] = imag_h_hold3_r[i];
        q_output_w[i] = q_output_r[i];
        mul_output2_w[i] = mul_output2_r[i];
        mul_output_w[i] = mul_output_r[i];
        
    end
    for(i=0;i<8;i=i+1)begin
        square_w[i]= {square_r[i],10'd0};
    end
    
    cnt_w = cnt_r;
    o_r_w = o_r_r;
    o_y_hat_w = o_y_hat_r;
    o_rd_vld_w = o_rd_vld_r;
    o_last_data_w = o_last_data_r;

    // div_val_w = div_val_r;
    count_2_w = count_2_r;
    cnt_out_w = cnt_out_r;

    real_h_hold1_w = real_h_hold1_r;
    imag_h_hold1_w = imag_h_hold1_r;
    real_h_hold2_w[0] = real_h_hold2_r[0];
    imag_h_hold2_w[0] = imag_h_hold2_r[0];
    real_h_hold2_w[1] = real_h_hold2_r[1];
    imag_h_hold2_w[1] = imag_h_hold2_r[1];

    div_val_w = div_val_r;

    o_r_hold_w = o_r_hold_r;
    cnt_w = (cnt_r == 5'd19)?5'd0:(i_trig||count_2_r==2'd2)?cnt_r + 1:cnt_r;
    mul_add = 0;
    if(i_trig)begin
        
        if(cnt_r==5'd4||cnt_r==5'd9||cnt_r==5'd14 ||cnt_r==5'd19)begin
            imag_origin_y_hold_w[cnt_r[1:0]] = i_data[47:38];
            real_origin_y_hold_w[cnt_r[1:0]] = i_data[23:14];
        end
        else begin
            if(cnt_r<5'd4)begin
                if(cnt_r==5'd0)begin
                    imag_h_w[0][0] = i_data[47:36];
                    real_h_w[0][0] = i_data[23:12];
                end
                else if(cnt_r==5'd1)begin
                    imag_h_hold1_w = i_data[47:36];
                    real_h_hold1_w = i_data[23:12];
                end
                else if(cnt_r==5'd2)begin
                    imag_h_hold2_w[0] = i_data[47:36];
                    real_h_hold2_w[0] = i_data[23:12];
                end
                else begin
                    imag_h_hold3_w[0] = i_data[47:36];
                    real_h_hold3_w[0] = i_data[23:12];
                end

            end
            else if(cnt_r<5'd9)begin
                if(cnt_r==5'd5)begin
                    imag_h_w[1][0] = i_data[47:36];
                    real_h_w[1][0] = i_data[23:12];
                end
                else if(cnt_r==5'd6)begin
                    imag_h_w[1][1] = i_data[47:36];
                    real_h_w[1][1] = i_data[23:12];
                end
                else if(cnt_r==5'd7)begin
                    imag_h_hold2_w[1] = i_data[47:36];
                    real_h_hold2_w[1] = i_data[23:12];
                end
                else begin
                    imag_h_hold3_w[1] = i_data[47:36];
                    real_h_hold3_w[1] = i_data[23:12];
                end

            end
            else if(cnt_r<5'd14)begin
                if(cnt_r==5'd10)begin
                    imag_h_w[2][0] = i_data[47:36];
                    real_h_w[2][0] = i_data[23:12];
                end
                else if(cnt_r==5'd11)begin
                    imag_h_w[2][1] = i_data[47:36];
                    real_h_w[2][1] = i_data[23:12];
                end
                else if(cnt_r==5'd12)begin
                    imag_h_w[2][2] = i_data[47:36];
                    real_h_w[2][2] = i_data[23:12];
                end
                else begin
                    imag_h_hold3_w[2] = i_data[47:36];
                    real_h_hold3_w[2] = i_data[23:12];
                end
            end
            else if(cnt_r<5'd19)begin
                if(cnt_r==5'd15)begin
                    imag_h_w[3][0] = i_data[47:36];
                    real_h_w[3][0] = i_data[23:12];
                end
                else if(cnt_r==5'd16)begin
                    imag_h_w[3][1] = i_data[47:36];
                    real_h_w[3][1] = i_data[23:12];
                end
                else if(cnt_r==5'd17)begin
                    imag_h_w[3][2] = i_data[47:36];
                    real_h_w[3][2] = i_data[23:12];
                end
                else begin
                    imag_h_hold3_w[3] = i_data[47:36];
                    real_h_hold3_w[3] = i_data[23:12];
                end

            end
        end
    end

    
    case (cnt_r)
        5'd16:begin
            //2
            real_h_w[0][3] = h_result[0];//h4(3)
            real_h_w[1][3] = h_result[1];
            real_h_w[2][3] = h_result[2];
            real_h_w[3][3] = h_result[3];
            imag_h_w[0][3] = h_result[4];
            imag_h_w[1][3] = h_result[5];
            imag_h_w[2][3] = h_result[6];
            imag_h_w[3][3] = h_result[7];
            

            count_2_w = (count_2_r==2'd2)?2'd2:count_2_r+1;
            
            for(i=0;i<8;i=i+1)begin
                square_w[i] = mul8_result[i][21:0];
            end
        end
        5'd17:begin
            o_r_hold_w[19:0] = {1'b0,sqrt_val[21:3]};//r11
            
            // {imag_h_w[0][1],real_h_w[0][1]} = {imag_h_r[0][1],real_h_r[0][1]};
            // {imag_h_w[1][1],real_h_w[1][1]} = {imag_h_r[1][1],real_h_r[1][1]};
            // {imag_h_w[2][1],real_h_w[2][1]} = {imag_h_r[2][1],real_h_r[2][1]};
            // {imag_h_w[3][1],real_h_w[3][1]} = {imag_h_r[3][1],real_h_r[3][1]};
            div_val_w = div_val_wire;
            for(i=0;i<8;i=i+1)begin
                square_w[i] = mul8_result[i][21:0];
            end
            mul_add = ((square_r[0] + square_r[1]) + (square_r[2] + square_r[3])) + ((square_r[4] + square_r[5]) + (square_r[6] + square_r[7]));
        end
        5'd18:begin
            
            q_w[0] = {mul8_result[0][22],mul8_result[0][19:1],mul8_result[4][22],mul8_result[4][19:1]};//e1
            q_w[1] = {mul8_result[1][22],mul8_result[1][19:1],mul8_result[5][22],mul8_result[5][19:1]};
            q_w[2] = {mul8_result[2][22],mul8_result[2][19:1],mul8_result[6][22],mul8_result[6][19:1]};
            q_w[3] = {mul8_result[3][22],mul8_result[3][19:1],mul8_result[7][22],mul8_result[7][19:1]};
            
            //2
            o_r_w[319:300] = {1'b0,sqrt_val[21:3]};//r44

            div_val_w = div_val_wire;

            if(cnt_out_r == 4'd8)begin
                o_last_data_w = 1;
            end
            mul_add = ((square_r[0] + square_r[1]) + (square_r[2] + square_r[3])) + ((square_r[4] + square_r[5]) + (square_r[6] + square_r[7]));
        end
        5'd19:begin
            //2
            q4_w[0] = {mul8_result[0][22],mul8_result[0][19:1],mul8_result[4][22],mul8_result[4][19:1]};//e4
            q4_w[1] = {mul8_result[1][22],mul8_result[1][19:1],mul8_result[5][22],mul8_result[5][19:1]};
            q4_w[2] = {mul8_result[2][22],mul8_result[2][19:1],mul8_result[6][22],mul8_result[6][19:1]};
            q4_w[3] = {mul8_result[3][22],mul8_result[3][19:1],mul8_result[7][22],mul8_result[7][19:1]};
            for(i=0;i<4;i=i+1)begin
                mul_output_w[i] = mul_output_wire[i];
            end
            o_last_data_w = 0;
            
        end
        5'd0:begin
            o_r_hold_w[59:20] = mul_output_add;//r12
            
            imag_h_w[0][3] = imag_h_hold3_r[0];
            real_h_w[0][3] = real_h_hold3_r[0];
            imag_h_w[1][3] = imag_h_hold3_r[1];
            real_h_w[1][3] = real_h_hold3_r[1];
            imag_h_w[2][3] = imag_h_hold3_r[2];
            real_h_w[2][3] = real_h_hold3_r[2];
            imag_h_w[3][3] = imag_h_hold3_r[3];
            real_h_w[3][3] = real_h_hold3_r[3];
            
            for(i=0;i<4;i=i+1)begin
                imag_origin_y_w[i] = imag_origin_y_hold_r[i];
                real_origin_y_w[i] = real_origin_y_hold_r[i];
            end
            for(i=0;i<4;i=i+1)begin
                q_output_w[i] ={y_and_mul2_out_wire[i][31:16],4'd0,y_and_mul2_out_wire[i][15:0],4'd0};
                mul_output_w[i] = mul_output_wire[i];
            end
            
        end
        5'd1:begin
            // o_r_w[119:80] = mul_output_add;//r13
            o_r_hold_w[99:60] = mul_output_add;//r13
            //2
            o_y_hat_w[139:120] = y_h_real; 
            o_y_hat_w[159:140] = y_h_imag;//y4
            o_rd_vld_w = (count_2_r==2'd2)?1:0;
            
            for(i=0;i<4;i=i+1)begin
                // q_output_w[i] = q_output_wire[i];
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
                mul_output_w[i] = mul_output_wire[i];
            end
            
        end
        5'd2:begin
            o_r_w[219:180] = mul_output_add;//r14
            o_r_w[59:0] = o_r_hold_r[59:0];//r11 r12
            o_r_w[119:80] = o_r_hold_r[99:60];//r13

            real_h_w[0][1] = h_result[0];//h2(1)
            real_h_w[1][1] = h_result[1];
            real_h_w[2][1] = h_result[2];
            real_h_w[3][1] = h_result[3];
            imag_h_w[0][1] = h_result[4];
            imag_h_w[1][1] = h_result[5];
            imag_h_w[2][1] = h_result[6];
            imag_h_w[3][1] = h_result[7];

            

            //2
            o_rd_vld_w = 0;
            cnt_out_w = (o_rd_vld_r&&cnt_out_r==4'd9)?0:(o_rd_vld_r)?cnt_out_r+1:cnt_out_r;
            // if(o_last_data_r)begin
            //     cnt_w = 0;
            //     count_2_w = 0;
            //     o_last_data_w = 0;
            // end
            for(i=0;i<4;i=i+1)begin
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
            end

            
        end
        5'd3:begin

            real_h_w[0][2] = h_result[0];//h3(1)
            real_h_w[1][2] = h_result[1];
            real_h_w[2][2] = h_result[2];
            real_h_w[3][2] = h_result[3];
            imag_h_w[0][2] = h_result[4];
            imag_h_w[1][2] = h_result[5];
            imag_h_w[2][2] = h_result[6];
            imag_h_w[3][2] = h_result[7];
            for(i=0;i<4;i=i+1)begin
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
            end
            for(i=0;i<8;i=i+1)begin
                square_w[i] = mul8_result[i][21:0];
            end
            
            for(i=0;i<4;i=i+1)begin
                imag_origin_y_w[i] = imag_origin_y_hold_r[i];
                real_origin_y_w[i] = real_origin_y_hold_r[i];
            end
        end
        5'd4:begin

            real_h_w[0][3] = h_result[0];//h4(1)
            real_h_w[1][3] = h_result[1];
            real_h_w[2][3] = h_result[2];
            real_h_w[3][3] = h_result[3];
            imag_h_w[0][3] = h_result[4];
            imag_h_w[1][3] = h_result[5];
            imag_h_w[2][3] = h_result[6];
            imag_h_w[3][3] = h_result[7];

            o_r_w[79:60] = {1'b0,sqrt_val[21:3]};//r22

            div_val_w = div_val_wire;

            for(i=0;i<4;i=i+1)begin
                q_output_w[i] ={y_and_mul2_out_wire[i][31:16],4'd0,y_and_mul2_out_wire[i][15:0],4'd0};
            end
            mul_add = ((square_r[0] + square_r[1]) + (square_r[2] + square_r[3])) + ((square_r[4] + square_r[5]) + (square_r[6] + square_r[7]));
        end
        5'd5:begin

            q_w[0] = {mul8_result[0][22],mul8_result[0][19:1],mul8_result[4][22],mul8_result[4][19:1]};//e2
            q_w[1] = {mul8_result[1][22],mul8_result[1][19:1],mul8_result[5][22],mul8_result[5][19:1]};
            q_w[2] = {mul8_result[2][22],mul8_result[2][19:1],mul8_result[6][22],mul8_result[6][19:1]};
            q_w[3] = {mul8_result[3][22],mul8_result[3][19:1],mul8_result[7][22],mul8_result[7][19:1]};

            o_y_hat_w[19:0] = y_h_real; 
            o_y_hat_w[39:20] = y_h_imag;//y1
        end
        5'd6:begin
            imag_h_w[0][1] = imag_h_hold1_r;
            real_h_w[0][1] = real_h_hold1_r;
            for(i=0;i<4;i=i+1)begin
                q_output_w[i] ={y_and_mul2_out_wire[i][31:16],4'd0,y_and_mul2_out_wire[i][15:0],4'd0};
                mul_output_w[i] = mul_output_wire[i];
            end
            
        end
        5'd7:begin
            o_r_w[159:120] = mul_output_add;//r23

            o_y_hat_w[59:40] = y_h_real; 
            o_y_hat_w[79:60] = y_h_imag;//y2
            for(i=0;i<4;i=i+1)begin
                mul_output_w[i] = mul_output_wire[i];
            end
        end
        5'd8:begin
            o_r_w[259:220] = mul_output_add;
            for(i=0;i<4;i=i+1)begin
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
            end
        end
        5'd9:begin
            real_h_w[0][2] = h_result[0];//h3(2)
            real_h_w[1][2] = h_result[1];
            real_h_w[2][2] = h_result[2];
            real_h_w[3][2] = h_result[3];
            imag_h_w[0][2] = h_result[4];
            imag_h_w[1][2] = h_result[5];
            imag_h_w[2][2] = h_result[6];
            imag_h_w[3][2] = h_result[7];

            for(i=0;i<4;i=i+1)begin
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
            end
        end
        5'd10:begin
            real_h_w[0][3] = h_result[0];//h4(2)
            real_h_w[1][3] = h_result[1];
            real_h_w[2][3] = h_result[2];
            real_h_w[3][3] = h_result[3];
            imag_h_w[0][3] = h_result[4];
            imag_h_w[1][3] = h_result[5];
            imag_h_w[2][3] = h_result[6];
            imag_h_w[3][3] = h_result[7];
            for(i=0;i<8;i=i+1)begin
                square_w[i] = mul8_result[i][21:0];
            end
        end
        5'd11:begin
            o_r_w[179:160] = {1'b0,sqrt_val[21:3]};//r33
            div_val_w = div_val_wire;
            mul_add = ((square_r[0] + square_r[1]) + (square_r[2] + square_r[3])) + ((square_r[4] + square_r[5]) + (square_r[6] + square_r[7]));
        end
        5'd12:begin

            q_w[0] = {mul8_result[0][22],mul8_result[0][19:1],mul8_result[4][22],mul8_result[4][19:1]};//e3
            q_w[1] = {mul8_result[1][22],mul8_result[1][19:1],mul8_result[5][22],mul8_result[5][19:1]};
            q_w[2] = {mul8_result[2][22],mul8_result[2][19:1],mul8_result[6][22],mul8_result[6][19:1]};
            q_w[3] = {mul8_result[3][22],mul8_result[3][19:1],mul8_result[7][22],mul8_result[7][19:1]};
        end
        5'd13:begin
            imag_h_w[0][2] = imag_h_hold2_r[0];
            real_h_w[0][2] = real_h_hold2_r[0];
            imag_h_w[1][2] = imag_h_hold2_r[1];
            real_h_w[1][2] = real_h_hold2_r[1];
            for(i=0;i<4;i=i+1)begin
                q_output_w[i] ={y_and_mul2_out_wire[i][31:16],4'd0,y_and_mul2_out_wire[i][15:0],4'd0};
                mul_output_w[i] = mul_output_wire[i];
            end
            
        end
        5'd14:begin
            o_r_w[299:260] = mul_output_add;


            
            o_y_hat_w[99:80] = y_h_real; 
            o_y_hat_w[119:100] = y_h_imag;//y3
            
        end
        5'd15:begin
            for(i=0;i<4;i=i+1)begin
                mul_output2_w[i] = {y_and_mul2_out_wire[i][31],y_and_mul2_out_wire[i][28:18],y_and_mul2_out_wire[i][15],y_and_mul2_out_wire[i][12:2]};
            end
        end
    endcase

end

always @(posedge i_clk or posedge i_rst) begin
    if(i_rst)begin
        for(i=0;i<4;i=i+1)begin
            for(j=0;j<4;j=j+1)begin
                real_h_r[i][j] <= 0;
                imag_h_r[i][j] <= 0;
                // real_h_hold_r[i][j] <= 0;
                // imag_h_hold_r[i][j] <= 0;
            end
            real_origin_y_r[i] <= 0;
            imag_origin_y_r[i] <= 0;
            q_r[i] <= 0;
            // q4_r[i] <= 0;

            mul_output_r[i] <= 0;
            mul_output2_r[i] <= 0;
            q_output_r[i] <= 0;
            imag_origin_y_hold_r[i] <= 0;
            real_origin_y_hold_r[i] <= 0;
            real_h_hold3_r[i] <= 0;
            imag_h_hold3_r[i] <= 0;
        end
        for(i=0;i<8;i=i+1)begin
            square_r[i]<= 0;
        end

        cnt_r <= 0;
        o_r_r <= 0;
        o_y_hat_r <= 0;
        o_rd_vld_r <= 0;
        o_last_data_r <= 0;

        div_val_r <= 0;
        count_2_r <= 0;
        cnt_out_r <= 0;
        
        o_r_hold_r <= 0;

        real_h_hold1_r <= 0;
        imag_h_hold1_r <= 0;
        real_h_hold2_r[0] <= 0;
        imag_h_hold2_r[0] <= 0;
        real_h_hold2_r[1] <= 0;
        imag_h_hold2_r[1] <= 0;
        
    end
    else begin
        for(i=0;i<4;i=i+1)begin
            for(j=0;j<4;j=j+1)begin
                real_h_r[i][j] <= real_h_w[i][j];
                imag_h_r[i][j] <= imag_h_w[i][j];
                // real_h_hold_r[i][j] <= real_h_hold_w[i][j];
                // imag_h_hold_r[i][j] <= imag_h_hold_w[i][j];
            end
            real_origin_y_r[i] <= real_origin_y_w[i];
            imag_origin_y_r[i] <= imag_origin_y_w[i];
            q_r[i] <= q_w[i];
            // q4_r[i] <= q4_w[i];

            mul_output_r[i] <= mul_output_w[i][39:0];
            mul_output2_r[i] <= mul_output2_w[i];
            q_output_r[i] <= (cnt_r ==5'd19)?q4_w[i]:q_output_w[i];
            imag_origin_y_hold_r[i] <= imag_origin_y_hold_w[i];
            real_origin_y_hold_r[i] <= real_origin_y_hold_w[i];
            real_h_hold3_r[i] <= real_h_hold3_w[i];
            imag_h_hold3_r[i] <= imag_h_hold3_w[i];
        end
        for(i=0;i<8;i=i+1)begin
            square_r[i]<= square_w[i][21:10];
        end

        cnt_r <= cnt_w;
        o_r_r <= o_r_w;
        o_y_hat_r <= o_y_hat_w;
        o_rd_vld_r <= o_rd_vld_w;
        o_last_data_r <= o_last_data_w;

        div_val_r <= div_val_w;
        count_2_r <= count_2_w;
        cnt_out_r <= cnt_out_w;
        o_r_hold_r <= o_r_hold_w;

        real_h_hold1_r <= real_h_hold1_w;
        imag_h_hold1_r <= imag_h_hold1_w;
        real_h_hold2_r[0] <= real_h_hold2_w[0];
        imag_h_hold2_r[0] <= imag_h_hold2_w[0];
        real_h_hold2_r[1] <= real_h_hold2_w[1];
        imag_h_hold2_r[1] <= imag_h_hold2_w[1];
    end
end
endmodule



module square_root_relate(
    input [14:0] sum,
    output reg [21:0] sqrt_val,
    output reg [21:0] div_val
);
    always @(*) begin
        case(sum[14:5])
            10'd0:begin
                sqrt_val = 22'b000_0010000000000000000;
                div_val= 22'b1000_000000000000000000;
            end
            10'd1:begin
                sqrt_val = 22'b000_0011011101101101000;
                div_val= 22'b0100_100111100110100111;
            end
            10'd2:begin
                sqrt_val = 22'b000_0100011110001101111;
                div_val= 22'b0011_100100111110010011;
            end
            10'd3:begin
                sqrt_val = 22'b000_0101010010101010000;
                div_val= 22'b0011_000001100001001001;
            end
            10'd4:begin
                sqrt_val = 22'b000_0110000000000000000;
                div_val= 22'b0010_101010101010101011;
            end
            10'd5:begin
                sqrt_val = 22'b000_0110101000100001110;
                div_val= 22'b0010_011010010111111011;
            end
            10'd6:begin
                sqrt_val = 22'b000_0111001101100000101;
                div_val= 22'b0010_001110000000001101;
            end
            10'd7:begin
                sqrt_val = 22'b000_0111101111101111100;
                div_val= 22'b0010_000100001100101010;
            end
            10'd8:begin
                sqrt_val = 22'b000_1000001111110000100;
                div_val= 22'b0001_111100001011011010;
            end
            10'd9:begin
                sqrt_val = 22'b000_1000101101111100001;
                div_val= 22'b0001_110101011101100000;
            end
            10'd10:begin
                sqrt_val = 22'b000_1001001010100100100;
                div_val= 22'b0001_101111101110100100;
            end
            10'd11:begin
                sqrt_val = 22'b000_1001100101110111100;
                div_val= 22'b0001_101010110000100110;
            end
            10'd12:begin
                sqrt_val = 22'b000_1010000000000000000;
                div_val= 22'b0001_100110011001100110;
            end
            10'd13:begin
                sqrt_val = 22'b000_1010011001000110111;
                div_val= 22'b0001_100010100010001101;
            end
            10'd14:begin
                sqrt_val = 22'b000_1010110001010011010;
                div_val= 22'b0001_011111000100110111;
            end
            10'd15:begin
                sqrt_val = 22'b000_1011001000101011001;
                div_val= 22'b0001_011011111101010100;
            end
            10'd16:begin
                sqrt_val = 22'b000_1011011111010011100;
                div_val= 22'b0001_011001001000001011;
            end
            10'd17:begin
                sqrt_val = 22'b000_1011110101010000100;
                div_val= 22'b0001_010110100010110011;
            end
            10'd18:begin
                sqrt_val = 22'b000_1100001010100110000;
                div_val= 22'b0001_010100001011000010;
            end
            10'd19:begin
                sqrt_val = 22'b000_1100011111010111000;
                div_val= 22'b0001_010001111111000101;
            end
            10'd20:begin
                sqrt_val = 22'b000_1100110011100110011;
                div_val= 22'b0001_001111111101100000;
            end
            10'd21:begin
                sqrt_val = 22'b000_1101000111010110100;
                div_val= 22'b0001_001110000101000101;
            end
            10'd22:begin
                sqrt_val = 22'b000_1101011010101001101;
                div_val= 22'b0001_001100010100110001;
            end
            10'd23:begin
                sqrt_val = 22'b000_1101101101100001100;
                div_val= 22'b0001_001010101011101101;
            end
            10'd24:begin
                sqrt_val = 22'b000_1110000000000000000;
                div_val= 22'b0001_001001001001001001;
            end
            10'd25:begin
                sqrt_val = 22'b000_1110010010000110101;
                div_val= 22'b0001_000111101100011100;
            end
            10'd26:begin
                sqrt_val = 22'b000_1110100011110110101;
                div_val= 22'b0001_000110010101000010;
            end
            10'd27:begin
                sqrt_val = 22'b000_1110110101010001100;
                div_val= 22'b0001_000101000010011100;
            end
            10'd28:begin
                sqrt_val = 22'b000_1111000110011000010;
                div_val= 22'b0001_000011110100001111;
            end
            10'd29:begin
                sqrt_val = 22'b000_1111010111001100000;
                div_val= 22'b0001_000010101010000010;
            end
            10'd30:begin
                sqrt_val = 22'b000_1111100111101101101;
                div_val= 22'b0001_000001100011100001;
            end
            10'd31:begin
                sqrt_val = 22'b000_1111110111111110000;
                div_val= 22'b0001_000000100000011000;
            end
            10'd32:begin
                sqrt_val = 22'b001_0000000111111110000;
                div_val= 22'b0000_111111100000011000;
            end
            10'd33:begin
                sqrt_val = 22'b001_0000010111101110011;
                div_val= 22'b0000_111110100011010000;
            end
            10'd34:begin
                sqrt_val = 22'b001_0000100111001111111;
                div_val= 22'b0000_111101101000110011;
            end
            10'd35:begin
                sqrt_val = 22'b001_0000110110100011000;
                div_val= 22'b0000_111100110000110110;
            end
            10'd36:begin
                sqrt_val = 22'b001_0001000101101000100;
                div_val= 22'b0000_111011111011001101;
            end
            10'd37:begin
                sqrt_val = 22'b001_0001010100100000110;
                div_val= 22'b0000_111011000111101110;
            end
            10'd38:begin
                sqrt_val = 22'b001_0001100011001100100;
                div_val= 22'b0000_111010010110010001;
            end
            10'd39:begin
                sqrt_val = 22'b001_0001110001101100001;
                div_val= 22'b0000_111001100110101100;
            end
            10'd40:begin
                sqrt_val = 22'b001_0010000000000000000;
                div_val= 22'b0000_111000111000111001;
            end
            10'd41:begin
                sqrt_val = 22'b001_0010001110001000101;
                div_val= 22'b0000_111000001100110000;
            end
            10'd42:begin
                sqrt_val = 22'b001_0010011100000110100;
                div_val= 22'b0000_110111100010001100;
            end
            10'd43:begin
                sqrt_val = 22'b001_0010101001111001111;
                div_val= 22'b0000_110110111001000110;
            end
            10'd44:begin
                sqrt_val = 22'b001_0010110111100011001;
                div_val= 22'b0000_110110010001011010;
            end
            10'd45:begin
                sqrt_val = 22'b001_0011000101000010110;
                div_val= 22'b0000_110101101011000001;
            end
            10'd46:begin
                sqrt_val = 22'b001_0011010010011000110;
                div_val= 22'b0000_110101000101111001;
            end
            10'd47:begin
                sqrt_val = 22'b001_0011011111100101110;
                div_val= 22'b0000_110100100001111011;
            end
            10'd48:begin
                sqrt_val = 22'b001_0011101100101001111;
                div_val= 22'b0000_110011111111000110;
            end
            10'd49:begin
                sqrt_val = 22'b001_0011111001100101011;
                div_val= 22'b0000_110011011101010100;
            end
            10'd50:begin
                sqrt_val = 22'b001_0100000110011000101;
                div_val= 22'b0000_110010111100100010;
            end
            10'd51:begin
                sqrt_val = 22'b001_0100010011000011110;
                div_val= 22'b0000_110010011100101111;
            end
            10'd52:begin
                sqrt_val = 22'b001_0100011111100111000;
                div_val= 22'b0000_110001111101110101;
            end
            10'd53:begin
                sqrt_val = 22'b001_0100101100000010110;
                div_val= 22'b0000_110001011111110011;
            end
            10'd54:begin
                sqrt_val = 22'b001_0100111000010111000;
                div_val= 22'b0000_110001000010100111;
            end
            10'd55:begin
                sqrt_val = 22'b001_0101000100100100001;
                div_val= 22'b0000_110000100110001101;
            end
            10'd56:begin
                sqrt_val = 22'b001_0101010000101010001;
                div_val= 22'b0000_110000001010100011;
            end
            10'd57:begin
                sqrt_val = 22'b001_0101011100101001011;
                div_val= 22'b0000_101111101111101000;
            end
            10'd58:begin
                sqrt_val = 22'b001_0101101000100010000;
                div_val= 22'b0000_101111010101011010;
            end
            10'd59:begin
                sqrt_val = 22'b001_0101110100010100001;
                div_val= 22'b0000_101110111011110110;
            end
            10'd60:begin
                sqrt_val = 22'b001_0110000000000000000;
                div_val= 22'b0000_101110100010111010;
            end
            10'd61:begin
                sqrt_val = 22'b001_0110001011100101101;
                div_val= 22'b0000_101110001010100110;
            end
            10'd62:begin
                sqrt_val = 22'b001_0110010111000101011;
                div_val= 22'b0000_101101110010110111;
            end
            10'd63:begin
                sqrt_val = 22'b001_0110100010011111001;
                div_val= 22'b0000_101101011011101100;
            end
            10'd64:begin
                sqrt_val = 22'b001_0110101101110011010;
                div_val= 22'b0000_101101000101000100;
            end
            10'd65:begin
                sqrt_val = 22'b001_0110111001000001110;
                div_val= 22'b0000_101100101110111101;
            end
            10'd66:begin
                sqrt_val = 22'b001_0111000100001010110;
                div_val= 22'b0000_101100011001010110;
            end
            10'd67:begin
                sqrt_val = 22'b001_0111001111001110100;
                div_val= 22'b0000_101100000100001110;
            end
            10'd68:begin
                sqrt_val = 22'b001_0111011010001100111;
                div_val= 22'b0000_101011101111100100;
            end
            10'd69:begin
                sqrt_val = 22'b001_0111100101000110010;
                div_val= 22'b0000_101011011011010110;
            end
            10'd70:begin
                sqrt_val = 22'b001_0111101111111010101;
                div_val= 22'b0000_101011000111100100;
            end
            10'd71:begin
                sqrt_val = 22'b001_0111111010101010001;
                div_val= 22'b0000_101010110100001101;
            end
            10'd72:begin
                sqrt_val = 22'b001_1000000101010100110;
                div_val= 22'b0000_101010100001001111;
            end
            10'd73:begin
                sqrt_val = 22'b001_1000001111111010110;
                div_val= 22'b0000_101010001110101010;
            end
            10'd74:begin
                sqrt_val = 22'b001_1000011010011100001;
                div_val= 22'b0000_101001111100011101;
            end
            10'd75:begin
                sqrt_val = 22'b001_1000100100111001000;
                div_val= 22'b0000_101001101010101000;
            end
            10'd76:begin
                sqrt_val = 22'b001_1000101111010001100;
                div_val= 22'b0000_101001011001001001;
            end
            10'd77:begin
                sqrt_val = 22'b001_1000111001100101101;
                div_val= 22'b0000_101001000111111111;
            end
            10'd78:begin
                sqrt_val = 22'b001_1001000011110101100;
                div_val= 22'b0000_101000110111001011;
            end
            10'd79:begin
                sqrt_val = 22'b001_1001001110000001010;
                div_val= 22'b0000_101000100110101011;
            end
            10'd80:begin
                sqrt_val = 22'b001_1001011000001000111;
                div_val= 22'b0000_101000010110011111;
            end
            10'd81:begin
                sqrt_val = 22'b001_1001100010001100100;
                div_val= 22'b0000_101000000110100110;
            end
            10'd82:begin
                sqrt_val = 22'b001_1001101100001100001;
                div_val= 22'b0000_100111110110111111;
            end
            10'd83:begin
                sqrt_val = 22'b001_1001110110001000000;
                div_val= 22'b0000_100111100111101010;
            end
            10'd84:begin
                sqrt_val = 22'b001_1010000000000000000;
                div_val= 22'b0000_100111011000100111;
            end
            10'd85:begin
                sqrt_val = 22'b001_1010001001110100010;
                div_val= 22'b0000_100111001001110101;
            end
            10'd86:begin
                sqrt_val = 22'b001_1010010011100100111;
                div_val= 22'b0000_100110111011010100;
            end
            10'd87:begin
                sqrt_val = 22'b001_1010011101010010000;
                div_val= 22'b0000_100110101101000010;
            end
            10'd88:begin
                sqrt_val = 22'b001_1010100110111011100;
                div_val= 22'b0000_100110011111000000;
            end
            10'd89:begin
                sqrt_val = 22'b001_1010110000100001100;
                div_val= 22'b0000_100110010001001100;
            end
            10'd90:begin
                sqrt_val = 22'b001_1010111010000100001;
                div_val= 22'b0000_100110000011101000;
            end
            10'd91:begin
                sqrt_val = 22'b001_1011000011100011011;
                div_val= 22'b0000_100101110110010010;
            end
            10'd92:begin
                sqrt_val = 22'b001_1011001100111111010;
                div_val= 22'b0000_100101101001001010;
            end
            10'd93:begin
                sqrt_val = 22'b001_1011010110010111111;
                div_val= 22'b0000_100101011100001111;
            end
            10'd94:begin
                sqrt_val = 22'b001_1011011111101101011;
                div_val= 22'b0000_100101001111100001;
            end
            10'd95:begin
                sqrt_val = 22'b001_1011101000111111110;
                div_val= 22'b0000_100101000011000001;
            end
            10'd96:begin
                sqrt_val = 22'b001_1011110010001110111;
                div_val= 22'b0000_100100110110101100;
            end
            10'd97:begin
                sqrt_val = 22'b001_1011111011011011000;
                div_val= 22'b0000_100100101010100100;
            end
            10'd98:begin
                sqrt_val = 22'b001_1100000100100100010;
                div_val= 22'b0000_100100011110101000;
            end
            10'd99:begin
                sqrt_val = 22'b001_1100001101101010011;
                div_val= 22'b0000_100100010010110111;
            end
            10'd100:begin
                sqrt_val = 22'b001_1100010110101101101;
                div_val= 22'b0000_100100000111010010;
            end
            10'd101:begin
                sqrt_val = 22'b001_1100011111101110000;
                div_val= 22'b0000_100011111011110111;
            end
            10'd102:begin
                sqrt_val = 22'b001_1100101000101011101;
                div_val= 22'b0000_100011110000100111;
            end
            10'd103:begin
                sqrt_val = 22'b001_1100110001100110011;
                div_val= 22'b0000_100011100101100010;
            end
            10'd104:begin
                sqrt_val = 22'b001_1100111010011110011;
                div_val= 22'b0000_100011011010100111;
            end
            10'd105:begin
                sqrt_val = 22'b001_1101000011010011101;
                div_val= 22'b0000_100011001111110110;
            end
            10'd106:begin
                sqrt_val = 22'b001_1101001100000110010;
                div_val= 22'b0000_100011000101001110;
            end
            10'd107:begin
                sqrt_val = 22'b001_1101010100110110010;
                div_val= 22'b0000_100010111010110001;
            end
            10'd108:begin
                sqrt_val = 22'b001_1101011101100011110;
                div_val= 22'b0000_100010110000011100;
            end
            10'd109:begin
                sqrt_val = 22'b001_1101100110001110100;
                div_val= 22'b0000_100010100110010000;
            end
            10'd110:begin
                sqrt_val = 22'b001_1101101110110110111;
                div_val= 22'b0000_100010011100001110;
            end
            10'd111:begin
                sqrt_val = 22'b001_1101110111011100101;
                div_val= 22'b0000_100010010010010100;
            end
            10'd112:begin
                sqrt_val = 22'b001_1110000000000000000;
                div_val= 22'b0000_100010001000100010;
            end
            10'd113:begin
                sqrt_val = 22'b001_1110001000100000111;
                div_val= 22'b0000_100001111110111001;
            end
            10'd114:begin
                sqrt_val = 22'b001_1110010000111111100;
                div_val= 22'b0000_100001110101011000;
            end
            10'd115:begin
                sqrt_val = 22'b001_1110011001011011101;
                div_val= 22'b0000_100001101011111110;
            end
            10'd116:begin
                sqrt_val = 22'b001_1110100001110101100;
                div_val= 22'b0000_100001100010101101;
            end
            10'd117:begin
                sqrt_val = 22'b001_1110101010001101000;
                div_val= 22'b0000_100001011001100011;
            end
            10'd118:begin
                sqrt_val = 22'b001_1110110010100010010;
                div_val= 22'b0000_100001010000100001;
            end
            10'd119:begin
                sqrt_val = 22'b001_1110111010110101010;
                div_val= 22'b0000_100001000111100101;
            end
            10'd120:begin
                sqrt_val = 22'b001_1111000011000110000;
                div_val= 22'b0000_100000111110110001;
            end
            10'd121:begin
                sqrt_val = 22'b001_1111001011010100101;
                div_val= 22'b0000_100000110110000100;
            end
            10'd122:begin
                sqrt_val = 22'b001_1111010011100001001;
                div_val= 22'b0000_100000101101011110;
            end
            10'd123:begin
                sqrt_val = 22'b001_1111011011101011011;
                div_val= 22'b0000_100000100100111111;
            end
            10'd124:begin
                sqrt_val = 22'b001_1111100011110011101;
                div_val= 22'b0000_100000011100100110;
            end
            10'd125:begin
                sqrt_val = 22'b001_1111101011111001110;
                div_val= 22'b0000_100000010100010011;
            end
            10'd126:begin
                sqrt_val = 22'b001_1111110011111101110;
                div_val= 22'b0000_100000001100000111;
            end
            10'd127:begin
                sqrt_val = 22'b001_1111111011111111110;
                div_val= 22'b0000_100000000100000001;
            end
            10'd128:begin
                sqrt_val = 22'b010_0000000011111111110;
                div_val= 22'b0000_011111111100000001;
            end
            10'd129:begin
                sqrt_val = 22'b010_0000001011111101110;
                div_val= 22'b0000_011111110100000111;
            end
            10'd130:begin
                sqrt_val = 22'b010_0000010011111001110;
                div_val= 22'b0000_011111101100010010;
            end
            10'd131:begin
                sqrt_val = 22'b010_0000011011110011111;
                div_val= 22'b0000_011111100100100100;
            end
            10'd132:begin
                sqrt_val = 22'b010_0000100011101100001;
                div_val= 22'b0000_011111011100111011;
            end
            10'd133:begin
                sqrt_val = 22'b010_0000101011100010011;
                div_val= 22'b0000_011111010101011000;
            end
            10'd134:begin
                sqrt_val = 22'b010_0000110011010110110;
                div_val= 22'b0000_011111001101111010;
            end
            10'd135:begin
                sqrt_val = 22'b010_0000111011001001011;
                div_val= 22'b0000_011111000110100001;
            end
            10'd136:begin
                sqrt_val = 22'b010_0001000010111010000;
                div_val= 22'b0000_011110111111001101;
            end
            10'd137:begin
                sqrt_val = 22'b010_0001001010101001000;
                div_val= 22'b0000_011110110111111111;
            end
            10'd138:begin
                sqrt_val = 22'b010_0001010010010110000;
                div_val= 22'b0000_011110110000110110;
            end
            10'd139:begin
                sqrt_val = 22'b010_0001011010000001011;
                div_val= 22'b0000_011110101001110001;
            end
            10'd140:begin
                sqrt_val = 22'b010_0001100001101011000;
                div_val= 22'b0000_011110100010110010;
            end
            10'd141:begin
                sqrt_val = 22'b010_0001101001010010110;
                div_val= 22'b0000_011110011011110111;
            end
            10'd142:begin
                sqrt_val = 22'b010_0001110000111000111;
                div_val= 22'b0000_011110010101000001;
            end
            10'd143:begin
                sqrt_val = 22'b010_0001111000011101010;
                div_val= 22'b0000_011110001110001111;
            end
            10'd144:begin
                sqrt_val = 22'b010_0010000000000000000;
                div_val= 22'b0000_011110000111100010;
            end
            10'd145:begin
                sqrt_val = 22'b010_0010000111100001000;
                div_val= 22'b0000_011110000000111001;
            end
            10'd146:begin
                sqrt_val = 22'b010_0010001111000000100;
                div_val= 22'b0000_011101111010010101;
            end
            10'd147:begin
                sqrt_val = 22'b010_0010010110011110010;
                div_val= 22'b0000_011101110011110101;
            end
            10'd148:begin
                sqrt_val = 22'b010_0010011101111010011;
                div_val= 22'b0000_011101101101011001;
            end
            10'd149:begin
                sqrt_val = 22'b010_0010100101010100111;
                div_val= 22'b0000_011101100111000001;
            end
            10'd150:begin
                sqrt_val = 22'b010_0010101100101101111;
                div_val= 22'b0000_011101100000101110;
            end
            10'd151:begin
                sqrt_val = 22'b010_0010110100000101010;
                div_val= 22'b0000_011101011010011110;
            end
            10'd152:begin
                sqrt_val = 22'b010_0010111011011011001;
                div_val= 22'b0000_011101010100010011;
            end
            10'd153:begin
                sqrt_val = 22'b010_0011000010101111011;
                div_val= 22'b0000_011101001110001011;
            end
            10'd154:begin
                sqrt_val = 22'b010_0011001010000010010;
                div_val= 22'b0000_011101001000000111;
            end
            10'd155:begin
                sqrt_val = 22'b010_0011010001010011100;
                div_val= 22'b0000_011101000010000111;
            end
            10'd156:begin
                sqrt_val = 22'b010_0011011000100011010;
                div_val= 22'b0000_011100111100001010;
            end
            10'd157:begin
                sqrt_val = 22'b010_0011011111110001101;
                div_val= 22'b0000_011100110110010001;
            end
            10'd158:begin
                sqrt_val = 22'b010_0011100110111110011;
                div_val= 22'b0000_011100110000011100;
            end
            10'd159:begin
                sqrt_val = 22'b010_0011101110001001110;
                div_val= 22'b0000_011100101010101010;
            end
            10'd160:begin
                sqrt_val = 22'b010_0011110101010011110;
                div_val= 22'b0000_011100100100111100;
            end
            10'd161:begin
                sqrt_val = 22'b010_0011111100011100010;
                div_val= 22'b0000_011100011111010001;
            end
            10'd162:begin
                sqrt_val = 22'b010_0100000011100011011;
                div_val= 22'b0000_011100011001101001;
            end
            10'd163:begin
                sqrt_val = 22'b010_0100001010101001001;
                div_val= 22'b0000_011100010100000101;
            end
            10'd164:begin
                sqrt_val = 22'b010_0100010001101101011;
                div_val= 22'b0000_011100001110100100;
            end
            10'd165:begin
                sqrt_val = 22'b010_0100011000110000011;
                div_val= 22'b0000_011100001001000110;
            end
            10'd166:begin
                sqrt_val = 22'b010_0100011111110010000;
                div_val= 22'b0000_011100000011101011;
            end
            10'd167:begin
                sqrt_val = 22'b010_0100100110110010010;
                div_val= 22'b0000_011011111110010100;
            end
            10'd168:begin
                sqrt_val = 22'b010_0100101101110001001;
                div_val= 22'b0000_011011111000111111;
            end
            10'd169:begin
                sqrt_val = 22'b010_0100110100101110110;
                div_val= 22'b0000_011011110011101110;
            end
            10'd170:begin
                sqrt_val = 22'b010_0100111011101011000;
                div_val= 22'b0000_011011101110011111;
            end
            10'd171:begin
                sqrt_val = 22'b010_0101000010100110000;
                div_val= 22'b0000_011011101001010100;
            end
            10'd172:begin
                sqrt_val = 22'b010_0101001001011111101;
                div_val= 22'b0000_011011100100001011;
            end
            10'd173:begin
                sqrt_val = 22'b010_0101010000011000000;
                div_val= 22'b0000_011011011111000101;
            end
            10'd174:begin
                sqrt_val = 22'b010_0101010111001111010;
                div_val= 22'b0000_011011011010000010;
            end
            10'd175:begin
                sqrt_val = 22'b010_0101011110000101001;
                div_val= 22'b0000_011011010101000010;
            end
            10'd176:begin
                sqrt_val = 22'b010_0101100100111001110;
                div_val= 22'b0000_011011010000000100;
            end
            10'd177:begin
                sqrt_val = 22'b010_0101101011101101001;
                div_val= 22'b0000_011011001011001001;
            end
            10'd178:begin
                sqrt_val = 22'b010_0101110010011111010;
                div_val= 22'b0000_011011000110010001;
            end
            10'd179:begin
                sqrt_val = 22'b010_0101111001010000010;
                div_val= 22'b0000_011011000001011011;
            end
            10'd180:begin
                sqrt_val = 22'b010_0110000000000000000;
                div_val= 22'b0000_011010111100101000;
            end
            10'd181:begin
                sqrt_val = 22'b010_0110000110101110100;
                div_val= 22'b0000_011010110111111000;
            end
            10'd182:begin
                sqrt_val = 22'b010_0110001101011100000;
                div_val= 22'b0000_011010110011001010;
            end
            10'd183:begin
                sqrt_val = 22'b010_0110010100001000001;
                div_val= 22'b0000_011010101110011110;
            end
            10'd184:begin
                sqrt_val = 22'b010_0110011010110011001;
                div_val= 22'b0000_011010101001110101;
            end
            10'd185:begin
                sqrt_val = 22'b010_0110100001011101001;
                div_val= 22'b0000_011010100101001111;
            end
            10'd186:begin
                sqrt_val = 22'b010_0110101000000101110;
                div_val= 22'b0000_011010100000101010;
            end
            10'd187:begin
                sqrt_val = 22'b010_0110101110101101011;
                div_val= 22'b0000_011010011100001000;
            end
            10'd188:begin
                sqrt_val = 22'b010_0110110101010011111;
                div_val= 22'b0000_011010010111101001;
            end
            10'd189:begin
                sqrt_val = 22'b010_0110111011111001010;
                div_val= 22'b0000_011010010011001011;
            end
            10'd190:begin
                sqrt_val = 22'b010_0111000010011101100;
                div_val= 22'b0000_011010001110110000;
            end
            10'd191:begin
                sqrt_val = 22'b010_0111001001000000101;
                div_val= 22'b0000_011010001010010111;
            end
            10'd192:begin
                sqrt_val = 22'b010_0111001111100010101;
                div_val= 22'b0000_011010000110000001;
            end
            10'd193:begin
                sqrt_val = 22'b010_0111010110000011101;
                div_val= 22'b0000_011010000001101100;
            end
            10'd194:begin
                sqrt_val = 22'b010_0111011100100011100;
                div_val= 22'b0000_011001111101011010;
            end
            10'd195:begin
                sqrt_val = 22'b010_0111100011000010011;
                div_val= 22'b0000_011001111001001010;
            end
            10'd196:begin
                sqrt_val = 22'b010_0111101001100000001;
                div_val= 22'b0000_011001110100111011;
            end
            10'd197:begin
                sqrt_val = 22'b010_0111101111111100110;
                div_val= 22'b0000_011001110000101111;
            end
            10'd198:begin
                sqrt_val = 22'b010_0111110110011000100;
                div_val= 22'b0000_011001101100100101;
            end
            10'd199:begin
                sqrt_val = 22'b010_0111111100110011001;
                div_val= 22'b0000_011001101000011101;
            end
            10'd200:begin
                sqrt_val = 22'b010_1000000011001100101;
                div_val= 22'b0000_011001100100010111;
            end
            10'd201:begin
                sqrt_val = 22'b010_1000001001100101010;
                div_val= 22'b0000_011001100000010011;
            end
            10'd202:begin
                sqrt_val = 22'b010_1000001111111100111;
                div_val= 22'b0000_011001011100010000;
            end
            10'd203:begin
                sqrt_val = 22'b010_1000010110010011011;
                div_val= 22'b0000_011001011000010000;
            end
            10'd204:begin
                sqrt_val = 22'b010_1000011100101001000;
                div_val= 22'b0000_011001010100010001;
            end
            10'd205:begin
                sqrt_val = 22'b010_1000100010111101100;
                div_val= 22'b0000_011001010000010101;
            end
            10'd206:begin
                sqrt_val = 22'b010_1000101001010001001;
                div_val= 22'b0000_011001001100011010;
            end
            10'd207:begin
                sqrt_val = 22'b010_1000101111100011110;
                div_val= 22'b0000_011001001000100001;
            end
            10'd208:begin
                sqrt_val = 22'b010_1000110101110101011;
                div_val= 22'b0000_011001000100101010;
            end
            10'd209:begin
                sqrt_val = 22'b010_1000111100000110000;
                div_val= 22'b0000_011001000000110101;
            end
            10'd210:begin
                sqrt_val = 22'b010_1001000010010101110;
                div_val= 22'b0000_011000111101000001;
            end
            10'd211:begin
                sqrt_val = 22'b010_1001001000100100101;
                div_val= 22'b0000_011000111001001111;
            end
            10'd212:begin
                sqrt_val = 22'b010_1001001110110010011;
                div_val= 22'b0000_011000110101011111;
            end
            10'd213:begin
                sqrt_val = 22'b010_1001010100111111010;
                div_val= 22'b0000_011000110001110000;
            end
            10'd214:begin
                sqrt_val = 22'b010_1001011011001011010;
                div_val= 22'b0000_011000101110000011;
            end
            10'd215:begin
                sqrt_val = 22'b010_1001100001010110011;
                div_val= 22'b0000_011000101010011000;
            end
            10'd216:begin
                sqrt_val = 22'b010_1001100111100000100;
                div_val= 22'b0000_011000100110101111;
            end
            10'd217:begin
                sqrt_val = 22'b010_1001101101101001110;
                div_val= 22'b0000_011000100011000111;
            end
            10'd218:begin
                sqrt_val = 22'b010_1001110011110010000;
                div_val= 22'b0000_011000011111100000;
            end
            10'd219:begin
                sqrt_val = 22'b010_1001111001111001100;
                div_val= 22'b0000_011000011011111100;
            end
            10'd220:begin
                sqrt_val = 22'b010_1010000000000000000;
                div_val= 22'b0000_011000011000011000;
            end
            10'd221:begin
                sqrt_val = 22'b010_1010000110000101101;
                div_val= 22'b0000_011000010100110111;
            end
            10'd222:begin
                sqrt_val = 22'b010_1010001100001010011;
                div_val= 22'b0000_011000010001010111;
            end
            10'd223:begin
                sqrt_val = 22'b010_1010010010001110011;
                div_val= 22'b0000_011000001101111000;
            end
            10'd224:begin
                sqrt_val = 22'b010_1010011000010001011;
                div_val= 22'b0000_011000001010011011;
            end
            10'd225:begin
                sqrt_val = 22'b010_1010011110010011100;
                div_val= 22'b0000_011000000110111111;
            end
            10'd226:begin
                sqrt_val = 22'b010_1010100100010100111;
                div_val= 22'b0000_011000000011100101;
            end
            10'd227:begin
                sqrt_val = 22'b010_1010101010010101011;
                div_val= 22'b0000_011000000000001100;
            end
            10'd228:begin
                sqrt_val = 22'b010_1010110000010101000;
                div_val= 22'b0000_010111111100110101;
            end
            10'd229:begin
                sqrt_val = 22'b010_1010110110010011110;
                div_val= 22'b0000_010111111001011111;
            end
            10'd230:begin
                sqrt_val = 22'b010_1010111100010001110;
                div_val= 22'b0000_010111110110001010;
            end
            10'd231:begin
                sqrt_val = 22'b010_1011000010001110111;
                div_val= 22'b0000_010111110010110111;
            end
            10'd232:begin
                sqrt_val = 22'b010_1011001000001011001;
                div_val= 22'b0000_010111101111100101;
            end
            10'd233:begin
                sqrt_val = 22'b010_1011001110000110101;
                div_val= 22'b0000_010111101100010101;
            end
            10'd234:begin
                sqrt_val = 22'b010_1011010100000001010;
                div_val= 22'b0000_010111101001000101;
            end
            10'd235:begin
                sqrt_val = 22'b010_1011011001111011001;
                div_val= 22'b0000_010111100101111000;
            end
            10'd236:begin
                sqrt_val = 22'b010_1011011111110100010;
                div_val= 22'b0000_010111100010101011;
            end
            10'd237:begin
                sqrt_val = 22'b010_1011100101101100100;
                div_val= 22'b0000_010111011111100000;
            end
            10'd238:begin
                sqrt_val = 22'b010_1011101011100100000;
                div_val= 22'b0000_010111011100010110;
            end
            10'd239:begin
                sqrt_val = 22'b010_1011110001011010101;
                div_val= 22'b0000_010111011001001101;
            end
            10'd240:begin
                sqrt_val = 22'b010_1011110111010000101;
                div_val= 22'b0000_010111010110000110;
            end
            10'd241:begin
                sqrt_val = 22'b010_1011111101000101110;
                div_val= 22'b0000_010111010011000000;
            end
            10'd242:begin
                sqrt_val = 22'b010_1100000010111010001;
                div_val= 22'b0000_010111001111111011;
            end
            10'd243:begin
                sqrt_val = 22'b010_1100001000101101101;
                div_val= 22'b0000_010111001100110111;
            end
            10'd244:begin
                sqrt_val = 22'b010_1100001110100000100;
                div_val= 22'b0000_010111001001110100;
            end
            10'd245:begin
                sqrt_val = 22'b010_1100010100010010101;
                div_val= 22'b0000_010111000110110011;
            end
            10'd246:begin
                sqrt_val = 22'b010_1100011010000011111;
                div_val= 22'b0000_010111000011110011;
            end
            10'd247:begin
                sqrt_val = 22'b010_1100011111110100100;
                div_val= 22'b0000_010111000000110100;
            end
            10'd248:begin
                sqrt_val = 22'b010_1100100101100100011;
                div_val= 22'b0000_010110111101110110;
            end
            10'd249:begin
                sqrt_val = 22'b010_1100101011010011011;
                div_val= 22'b0000_010110111010111001;
            end
            10'd250:begin
                sqrt_val = 22'b010_1100110001000001110;
                div_val= 22'b0000_010110110111111110;
            end
            10'd251:begin
                sqrt_val = 22'b010_1100110110101111011;
                div_val= 22'b0000_010110110101000011;
            end
            10'd252:begin
                sqrt_val = 22'b010_1100111100011100010;
                div_val= 22'b0000_010110110010001010;
            end
            10'd253:begin
                sqrt_val = 22'b010_1101000010001000100;
                div_val= 22'b0000_010110101111010010;
            end
            10'd254:begin
                sqrt_val = 22'b010_1101000111110100000;
                div_val= 22'b0000_010110101100011011;
            end
            10'd255:begin
                sqrt_val = 22'b010_1101001101011110110;
                div_val= 22'b0000_010110101001100101;
            end
            10'd256:begin
                sqrt_val = 22'b010_1101010011001000110;
                div_val= 22'b0000_010110100110110000;
            end
            10'd257:begin
                sqrt_val = 22'b010_1101011000110010001;
                div_val= 22'b0000_010110100011111100;
            end
            10'd258:begin
                sqrt_val = 22'b010_1101011110011010110;
                div_val= 22'b0000_010110100001001001;
            end
            10'd259:begin
                sqrt_val = 22'b010_1101100100000010101;
                div_val= 22'b0000_010110011110010111;
            end
            10'd260:begin
                sqrt_val = 22'b010_1101101001101001111;
                div_val= 22'b0000_010110011011100110;
            end
            10'd261:begin
                sqrt_val = 22'b010_1101101111010000011;
                div_val= 22'b0000_010110011000110110;
            end
            10'd262:begin
                sqrt_val = 22'b010_1101110100110110010;
                div_val= 22'b0000_010110010110000111;
            end
            10'd263:begin
                sqrt_val = 22'b010_1101111010011011100;
                div_val= 22'b0000_010110010011011001;
            end
            10'd264:begin
                sqrt_val = 22'b010_1110000000000000000;
                div_val= 22'b0000_010110010000101101;
            end
            10'd265:begin
                sqrt_val = 22'b010_1110000101100011111;
                div_val= 22'b0000_010110001110000001;
            end
            10'd266:begin
                sqrt_val = 22'b010_1110001011000111000;
                div_val= 22'b0000_010110001011010110;
            end
            10'd267:begin
                sqrt_val = 22'b010_1110010000101001100;
                div_val= 22'b0000_010110001000101100;
            end
            10'd268:begin
                sqrt_val = 22'b010_1110010110001011011;
                div_val= 22'b0000_010110000110000011;
            end
            10'd269:begin
                sqrt_val = 22'b010_1110011011101100100;
                div_val= 22'b0000_010110000011011011;
            end
            10'd270:begin
                sqrt_val = 22'b010_1110100001001101000;
                div_val= 22'b0000_010110000000110100;
            end
            10'd271:begin
                sqrt_val = 22'b010_1110100110101100111;
                div_val= 22'b0000_010101111110001101;
            end
            10'd272:begin
                sqrt_val = 22'b010_1110101100001100001;
                div_val= 22'b0000_010101111011101000;
            end
            10'd273:begin
                sqrt_val = 22'b010_1110110001101010110;
                div_val= 22'b0000_010101111001000100;
            end
            10'd274:begin
                sqrt_val = 22'b010_1110110111001000110;
                div_val= 22'b0000_010101110110100000;
            end
            10'd275:begin
                sqrt_val = 22'b010_1110111100100110000;
                div_val= 22'b0000_010101110011111110;
            end
            10'd276:begin
                sqrt_val = 22'b010_1111000010000010101;
                div_val= 22'b0000_010101110001011100;
            end
            10'd277:begin
                sqrt_val = 22'b010_1111000111011110110;
                div_val= 22'b0000_010101101110111011;
            end
            10'd278:begin
                sqrt_val = 22'b010_1111001100111010001;
                div_val= 22'b0000_010101101100011011;
            end
            10'd279:begin
                sqrt_val = 22'b010_1111010010010100111;
                div_val= 22'b0000_010101101001111100;
            end
            10'd280:begin
                sqrt_val = 22'b010_1111010111101111001;
                div_val= 22'b0000_010101100111011110;
            end
            10'd281:begin
                sqrt_val = 22'b010_1111011101001000101;
                div_val= 22'b0000_010101100101000000;
            end
            10'd282:begin
                sqrt_val = 22'b010_1111100010100001101;
                div_val= 22'b0000_010101100010100100;
            end
            10'd283:begin
                sqrt_val = 22'b010_1111100111111010000;
                div_val= 22'b0000_010101100000001000;
            end
            10'd284:begin
                sqrt_val = 22'b010_1111101101010001101;
                div_val= 22'b0000_010101011101101101;
            end
            10'd285:begin
                sqrt_val = 22'b010_1111110010101000110;
                div_val= 22'b0000_010101011011010011;
            end
            10'd286:begin
                sqrt_val = 22'b010_1111110111111111011;
                div_val= 22'b0000_010101011000111010;
            end
            10'd287:begin
                sqrt_val = 22'b010_1111111101010101010;
                div_val= 22'b0000_010101010110100001;
            end
            10'd288:begin
                sqrt_val = 22'b011_0000000010101010101;
                div_val= 22'b0000_010101010100001010;
            end
            10'd289:begin
                sqrt_val = 22'b011_0000000111111111011;
                div_val= 22'b0000_010101010001110011;
            end
            10'd290:begin
                sqrt_val = 22'b011_0000001101010011100;
                div_val= 22'b0000_010101001111011101;
            end
            10'd291:begin
                sqrt_val = 22'b011_0000010010100111000;
                div_val= 22'b0000_010101001101000111;
            end
            10'd292:begin
                sqrt_val = 22'b011_0000010111111010000;
                div_val= 22'b0000_010101001010110011;
            end
            10'd293:begin
                sqrt_val = 22'b011_0000011101001100100;
                div_val= 22'b0000_010101001000011111;
            end
            10'd294:begin
                sqrt_val = 22'b011_0000100010011110010;
                div_val= 22'b0000_010101000110001100;
            end
            10'd295:begin
                sqrt_val = 22'b011_0000100111101111100;
                div_val= 22'b0000_010101000011111001;
            end
            10'd296:begin
                sqrt_val = 22'b011_0000101101000000010;
                div_val= 22'b0000_010101000001101000;
            end
            10'd297:begin
                sqrt_val = 22'b011_0000110010010000011;
                div_val= 22'b0000_010100111111010111;
            end
            10'd298:begin
                sqrt_val = 22'b011_0000110111011111111;
                div_val= 22'b0000_010100111101000111;
            end
            10'd299:begin
                sqrt_val = 22'b011_0000111100101110111;
                div_val= 22'b0000_010100111010110111;
            end
            10'd300:begin
                sqrt_val = 22'b011_0001000001111101011;
                div_val= 22'b0000_010100111000101001;
            end
            10'd301:begin
                sqrt_val = 22'b011_0001000111001011010;
                div_val= 22'b0000_010100110110011011;
            end
            10'd302:begin
                sqrt_val = 22'b011_0001001100011000100;
                div_val= 22'b0000_010100110100001101;
            end
            10'd303:begin
                sqrt_val = 22'b011_0001010001100101011;
                div_val= 22'b0000_010100110010000001;
            end
            10'd304:begin
                sqrt_val = 22'b011_0001010110110001101;
                div_val= 22'b0000_010100101111110101;
            end
            10'd305:begin
                sqrt_val = 22'b011_0001011011111101010;
                div_val= 22'b0000_010100101101101010;
            end
            10'd306:begin
                sqrt_val = 22'b011_0001100001001000011;
                div_val= 22'b0000_010100101011011111;
            end
            10'd307:begin
                sqrt_val = 22'b011_0001100110010011000;
                div_val= 22'b0000_010100101001010101;
            end
            10'd308:begin
                sqrt_val = 22'b011_0001101011011101000;
                div_val= 22'b0000_010100100111001100;
            end
            10'd309:begin
                sqrt_val = 22'b011_0001110000100110101;
                div_val= 22'b0000_010100100101000100;
            end
            10'd310:begin
                sqrt_val = 22'b011_0001110101101111101;
                div_val= 22'b0000_010100100010111100;
            end
            10'd311:begin
                sqrt_val = 22'b011_0001111010111000000;
                div_val= 22'b0000_010100100000110101;
            end
            10'd312:begin
                sqrt_val = 22'b011_0010000000000000000;
                div_val= 22'b0000_010100011110101110;
            end
            10'd313:begin
                sqrt_val = 22'b011_0010000101000111011;
                div_val= 22'b0000_010100011100101000;
            end
            10'd314:begin
                sqrt_val = 22'b011_0010001010001110011;
                div_val= 22'b0000_010100011010100011;
            end
            10'd315:begin
                sqrt_val = 22'b011_0010001111010100110;
                div_val= 22'b0000_010100011000011110;
            end
            10'd316:begin
                sqrt_val = 22'b011_0010010100011010100;
                div_val= 22'b0000_010100010110011010;
            end
            10'd317:begin
                sqrt_val = 22'b011_0010011001011111111;
                div_val= 22'b0000_010100010100010111;
            end
            10'd318:begin
                sqrt_val = 22'b011_0010011110100100110;
                div_val= 22'b0000_010100010010010100;
            end
            10'd319:begin
                sqrt_val = 22'b011_0010100011101001000;
                div_val= 22'b0000_010100010000010010;
            end
            10'd320:begin
                sqrt_val = 22'b011_0010101000101100111;
                div_val= 22'b0000_010100001110010001;
            end
            10'd321:begin
                sqrt_val = 22'b011_0010101101110000001;
                div_val= 22'b0000_010100001100010000;
            end
            10'd322:begin
                sqrt_val = 22'b011_0010110010110011000;
                div_val= 22'b0000_010100001010001111;
            end
            10'd323:begin
                sqrt_val = 22'b011_0010110111110101010;
                div_val= 22'b0000_010100001000010000;
            end
            10'd324:begin
                sqrt_val = 22'b011_0010111100110111001;
                div_val= 22'b0000_010100000110010000;
            end
            10'd325:begin
                sqrt_val = 22'b011_0011000001111000011;
                div_val= 22'b0000_010100000100010010;
            end
            10'd326:begin
                sqrt_val = 22'b011_0011000110111001010;
                div_val= 22'b0000_010100000010010100;
            end
            10'd327:begin
                sqrt_val = 22'b011_0011001011111001101;
                div_val= 22'b0000_010100000000010111;
            end
            10'd328:begin
                sqrt_val = 22'b011_0011010000111001011;
                div_val= 22'b0000_010011111110011010;
            end
            10'd329:begin
                sqrt_val = 22'b011_0011010101111000110;
                div_val= 22'b0000_010011111100011101;
            end
            10'd330:begin
                sqrt_val = 22'b011_0011011010110111101;
                div_val= 22'b0000_010011111010100010;
            end
            10'd331:begin
                sqrt_val = 22'b011_0011011111110110000;
                div_val= 22'b0000_010011111000100111;
            end
            10'd332:begin
                sqrt_val = 22'b011_0011100100110100000;
                div_val= 22'b0000_010011110110101100;
            end
            10'd333:begin
                sqrt_val = 22'b011_0011101001110001011;
                div_val= 22'b0000_010011110100110010;
            end
            10'd334:begin
                sqrt_val = 22'b011_0011101110101110011;
                div_val= 22'b0000_010011110010111001;
            end
            10'd335:begin
                sqrt_val = 22'b011_0011110011101010111;
                div_val= 22'b0000_010011110001000000;
            end
            10'd336:begin
                sqrt_val = 22'b011_0011111000100110111;
                div_val= 22'b0000_010011101111000111;
            end
            10'd337:begin
                sqrt_val = 22'b011_0011111101100010011;
                div_val= 22'b0000_010011101101001111;
            end
            10'd338:begin
                sqrt_val = 22'b011_0100000010011101100;
                div_val= 22'b0000_010011101011011000;
            end
            10'd339:begin
                sqrt_val = 22'b011_0100000111011000001;
                div_val= 22'b0000_010011101001100001;
            end
            10'd340:begin
                sqrt_val = 22'b011_0100001100010010010;
                div_val= 22'b0000_010011100111101011;
            end
            10'd341:begin
                sqrt_val = 22'b011_0100010001001011111;
                div_val= 22'b0000_010011100101110101;
            end
            10'd342:begin
                sqrt_val = 22'b011_0100010110000101001;
                div_val= 22'b0000_010011100100000000;
            end
            10'd343:begin
                sqrt_val = 22'b011_0100011010111101111;
                div_val= 22'b0000_010011100010001011;
            end
            10'd344:begin
                sqrt_val = 22'b011_0100011111110110010;
                div_val= 22'b0000_010011100000010111;
            end
            10'd345:begin
                sqrt_val = 22'b011_0100100100101110001;
                div_val= 22'b0000_010011011110100011;
            end
            10'd346:begin
                sqrt_val = 22'b011_0100101001100101100;
                div_val= 22'b0000_010011011100110000;
            end
            10'd347:begin
                sqrt_val = 22'b011_0100101110011100100;
                div_val= 22'b0000_010011011010111110;
            end
            10'd348:begin
                sqrt_val = 22'b011_0100110011010011000;
                div_val= 22'b0000_010011011001001011;
            end
            10'd349:begin
                sqrt_val = 22'b011_0100111000001001001;
                div_val= 22'b0000_010011010111011010;
            end
            10'd350:begin
                sqrt_val = 22'b011_0100111100111110110;
                div_val= 22'b0000_010011010101101000;
            end
            10'd351:begin
                sqrt_val = 22'b011_0101000001110011111;
                div_val= 22'b0000_010011010011111000;
            end
            10'd352:begin
                sqrt_val = 22'b011_0101000110101000101;
                div_val= 22'b0000_010011010010000111;
            end
            10'd353:begin
                sqrt_val = 22'b011_0101001011011101000;
                div_val= 22'b0000_010011010000011000;
            end
            10'd354:begin
                sqrt_val = 22'b011_0101010000010000111;
                div_val= 22'b0000_010011001110101000;
            end
            10'd355:begin
                sqrt_val = 22'b011_0101010101000100010;
                div_val= 22'b0000_010011001100111001;
            end
            10'd356:begin
                sqrt_val = 22'b011_0101011001110111010;
                div_val= 22'b0000_010011001011001011;
            end
            10'd357:begin
                sqrt_val = 22'b011_0101011110101001111;
                div_val= 22'b0000_010011001001011101;
            end
            10'd358:begin
                sqrt_val = 22'b011_0101100011011100000;
                div_val= 22'b0000_010011000111110000;
            end
            10'd359:begin
                sqrt_val = 22'b011_0101101000001101110;
                div_val= 22'b0000_010011000110000011;
            end
            10'd360:begin
                sqrt_val = 22'b011_0101101100111111000;
                div_val= 22'b0000_010011000100010110;
            end
            10'd361:begin
                sqrt_val = 22'b011_0101110001101111111;
                div_val= 22'b0000_010011000010101010;
            end
            10'd362:begin
                sqrt_val = 22'b011_0101110110100000011;
                div_val= 22'b0000_010011000000111110;
            end
            10'd363:begin
                sqrt_val = 22'b011_0101111011010000011;
                div_val= 22'b0000_010010111111010011;
            end
            10'd364:begin
                sqrt_val = 22'b011_0110000000000000000;
                div_val= 22'b0000_010010111101101000;
            end
            10'd365:begin
                sqrt_val = 22'b011_0110000100101111010;
                div_val= 22'b0000_010010111011111110;
            end
            10'd366:begin
                sqrt_val = 22'b011_0110001001011110000;
                div_val= 22'b0000_010010111010010100;
            end
            10'd367:begin
                sqrt_val = 22'b011_0110001110001100011;
                div_val= 22'b0000_010010111000101011;
            end
            10'd368:begin
                sqrt_val = 22'b011_0110010010111010011;
                div_val= 22'b0000_010010110111000010;
            end
            10'd369:begin
                sqrt_val = 22'b011_0110010111100111111;
                div_val= 22'b0000_010010110101011001;
            end
            10'd370:begin
                sqrt_val = 22'b011_0110011100010101000;
                div_val= 22'b0000_010010110011110001;
            end
            10'd371:begin
                sqrt_val = 22'b011_0110100001000001110;
                div_val= 22'b0000_010010110010001001;
            end
            10'd372:begin
                sqrt_val = 22'b011_0110100101101110001;
                div_val= 22'b0000_010010110000100010;
            end
            10'd373:begin
                sqrt_val = 22'b011_0110101010011010000;
                div_val= 22'b0000_010010101110111011;
            end
            10'd374:begin
                sqrt_val = 22'b011_0110101111000101100;
                div_val= 22'b0000_010010101101010100;
            end
            10'd375:begin
                sqrt_val = 22'b011_0110110011110000101;
                div_val= 22'b0000_010010101011101110;
            end
            10'd376:begin
                sqrt_val = 22'b011_0110111000011011011;
                div_val= 22'b0000_010010101010001000;
            end
            10'd377:begin
                sqrt_val = 22'b011_0110111101000101110;
                div_val= 22'b0000_010010101000100011;
            end
            10'd378:begin
                sqrt_val = 22'b011_0111000001101111101;
                div_val= 22'b0000_010010100110111110;
            end
            10'd379:begin
                sqrt_val = 22'b011_0111000110011001010;
                div_val= 22'b0000_010010100101011010;
            end
            10'd380:begin
                sqrt_val = 22'b011_0111001011000010011;
                div_val= 22'b0000_010010100011110110;
            end
            10'd381:begin
                sqrt_val = 22'b011_0111001111101011001;
                div_val= 22'b0000_010010100010010010;
            end
            10'd382:begin
                sqrt_val = 22'b011_0111010100010011100;
                div_val= 22'b0000_010010100000101111;
            end
            10'd383:begin
                sqrt_val = 22'b011_0111011000111011100;
                div_val= 22'b0000_010010011111001100;
            end
            10'd384:begin
                sqrt_val = 22'b011_0111011101100011001;
                div_val= 22'b0000_010010011101101001;
            end
            10'd385:begin
                sqrt_val = 22'b011_0111100010001010011;
                div_val= 22'b0000_010010011100000111;
            end
            10'd386:begin
                sqrt_val = 22'b011_0111100110110001001;
                div_val= 22'b0000_010010011010100101;
            end
            10'd387:begin
                sqrt_val = 22'b011_0111101011010111101;
                div_val= 22'b0000_010010011001000100;
            end
            10'd388:begin
                sqrt_val = 22'b011_0111101111111101110;
                div_val= 22'b0000_010010010111100011;
            end
            10'd389:begin
                sqrt_val = 22'b011_0111110100100011011;
                div_val= 22'b0000_010010010110000010;
            end
            10'd390:begin
                sqrt_val = 22'b011_0111111001001000110;
                div_val= 22'b0000_010010010100100010;
            end
            10'd391:begin
                sqrt_val = 22'b011_0111111101101101101;
                div_val= 22'b0000_010010010011000010;
            end
            10'd392:begin
                sqrt_val = 22'b011_1000000010010010010;
                div_val= 22'b0000_010010010001100011;
            end
            10'd393:begin
                sqrt_val = 22'b011_1000000110110110100;
                div_val= 22'b0000_010010010000000011;
            end
            10'd394:begin
                sqrt_val = 22'b011_1000001011011010010;
                div_val= 22'b0000_010010001110100101;
            end
            10'd395:begin
                sqrt_val = 22'b011_1000001111111101110;
                div_val= 22'b0000_010010001101000110;
            end
            10'd396:begin
                sqrt_val = 22'b011_1000010100100000111;
                div_val= 22'b0000_010010001011101000;
            end
            10'd397:begin
                sqrt_val = 22'b011_1000011001000011100;
                div_val= 22'b0000_010010001010001010;
            end
            10'd398:begin
                sqrt_val = 22'b011_1000011101100101111;
                div_val= 22'b0000_010010001000101101;
            end
            10'd399:begin
                sqrt_val = 22'b011_1000100010000111111;
                div_val= 22'b0000_010010000111010000;
            end
            10'd400:begin
                sqrt_val = 22'b011_1000100110101001100;
                div_val= 22'b0000_010010000101110011;
            end
            10'd401:begin
                sqrt_val = 22'b011_1000101011001010110;
                div_val= 22'b0000_010010000100010111;
            end
            10'd402:begin
                sqrt_val = 22'b011_1000101111101011110;
                div_val= 22'b0000_010010000010111011;
            end
            10'd403:begin
                sqrt_val = 22'b011_1000110100001100010;
                div_val= 22'b0000_010010000001011111;
            end
            10'd404:begin
                sqrt_val = 22'b011_1000111000101100100;
                div_val= 22'b0000_010010000000000100;
            end
            10'd405:begin
                sqrt_val = 22'b011_1000111101001100010;
                div_val= 22'b0000_010001111110101001;
            end
            10'd406:begin
                sqrt_val = 22'b011_1001000001101011110;
                div_val= 22'b0000_010001111101001110;
            end
            10'd407:begin
                sqrt_val = 22'b011_1001000110001010111;
                div_val= 22'b0000_010001111011110100;
            end
            10'd408:begin
                sqrt_val = 22'b011_1001001010101001101;
                div_val= 22'b0000_010001111010011010;
            end
            10'd409:begin
                sqrt_val = 22'b011_1001001111001000001;
                div_val= 22'b0000_010001111001000000;
            end
            10'd410:begin
                sqrt_val = 22'b011_1001010011100110001;
                div_val= 22'b0000_010001110111100111;
            end
            10'd411:begin
                sqrt_val = 22'b011_1001011000000011111;
                div_val= 22'b0000_010001110110001110;
            end
            10'd412:begin
                sqrt_val = 22'b011_1001011100100001010;
                div_val= 22'b0000_010001110100110101;
            end
            10'd413:begin
                sqrt_val = 22'b011_1001100000111110011;
                div_val= 22'b0000_010001110011011101;
            end
            10'd414:begin
                sqrt_val = 22'b011_1001100101011011000;
                div_val= 22'b0000_010001110010000101;
            end
            10'd415:begin
                sqrt_val = 22'b011_1001101001110111011;
                div_val= 22'b0000_010001110000101101;
            end
            10'd416:begin
                sqrt_val = 22'b011_1001101110010011011;
                div_val= 22'b0000_010001101111010110;
            end
            10'd417:begin
                sqrt_val = 22'b011_1001110010101111000;
                div_val= 22'b0000_010001101101111111;
            end
            10'd418:begin
                sqrt_val = 22'b011_1001110111001010011;
                div_val= 22'b0000_010001101100101000;
            end
            10'd419:begin
                sqrt_val = 22'b011_1001111011100101011;
                div_val= 22'b0000_010001101011010010;
            end
            10'd420:begin
                sqrt_val = 22'b011_1010000000000000000;
                div_val= 22'b0000_010001101001111100;
            end
            10'd421:begin
                sqrt_val = 22'b011_1010000100011010011;
                div_val= 22'b0000_010001101000100110;
            end
            10'd422:begin
                sqrt_val = 22'b011_1010001000110100010;
                div_val= 22'b0000_010001100111010000;
            end
            10'd423:begin
                sqrt_val = 22'b011_1010001101001110000;
                div_val= 22'b0000_010001100101111011;
            end
            10'd424:begin
                sqrt_val = 22'b011_1010010001100111010;
                div_val= 22'b0000_010001100100100110;
            end
            10'd425:begin
                sqrt_val = 22'b011_1010010110000000010;
                div_val= 22'b0000_010001100011010001;
            end
            10'd426:begin
                sqrt_val = 22'b011_1010011010011000111;
                div_val= 22'b0000_010001100001111101;
            end
            10'd427:begin
                sqrt_val = 22'b011_1010011110110001010;
                div_val= 22'b0000_010001100000101001;
            end
            10'd428:begin
                sqrt_val = 22'b011_1010100011001001010;
                div_val= 22'b0000_010001011111010101;
            end
            10'd429:begin
                sqrt_val = 22'b011_1010100111100000111;
                div_val= 22'b0000_010001011110000010;
            end
            10'd430:begin
                sqrt_val = 22'b011_1010101011111000010;
                div_val= 22'b0000_010001011100101111;
            end
            10'd431:begin
                sqrt_val = 22'b011_1010110000001111010;
                div_val= 22'b0000_010001011011011100;
            end
            10'd432:begin
                sqrt_val = 22'b011_1010110100100110000;
                div_val= 22'b0000_010001011010001001;
            end
            10'd433:begin
                sqrt_val = 22'b011_1010111000111100011;
                div_val= 22'b0000_010001011000110111;
            end
            10'd434:begin
                sqrt_val = 22'b011_1010111101010010011;
                div_val= 22'b0000_010001010111100101;
            end
            10'd435:begin
                sqrt_val = 22'b011_1011000001101000001;
                div_val= 22'b0000_010001010110010011;
            end
            10'd436:begin
                sqrt_val = 22'b011_1011000101111101100;
                div_val= 22'b0000_010001010101000010;
            end
            10'd437:begin
                sqrt_val = 22'b011_1011001010010010101;
                div_val= 22'b0000_010001010011110001;
            end
            10'd438:begin
                sqrt_val = 22'b011_1011001110100111011;
                div_val= 22'b0000_010001010010100000;
            end
            10'd439:begin
                sqrt_val = 22'b011_1011010010111011111;
                div_val= 22'b0000_010001010001001111;
            end
            10'd440:begin
                sqrt_val = 22'b011_1011010111010000000;
                div_val= 22'b0000_010001001111111111;
            end
            10'd441:begin
                sqrt_val = 22'b011_1011011011100011111;
                div_val= 22'b0000_010001001110101111;
            end
            10'd442:begin
                sqrt_val = 22'b011_1011011111110111011;
                div_val= 22'b0000_010001001101011111;
            end
            10'd443:begin
                sqrt_val = 22'b011_1011100100001010101;
                div_val= 22'b0000_010001001100001111;
            end
            10'd444:begin
                sqrt_val = 22'b011_1011101000011101100;
                div_val= 22'b0000_010001001011000000;
            end
            10'd445:begin
                sqrt_val = 22'b011_1011101100110000001;
                div_val= 22'b0000_010001001001110001;
            end
            10'd446:begin
                sqrt_val = 22'b011_1011110001000010011;
                div_val= 22'b0000_010001001000100011;
            end
            10'd447:begin
                sqrt_val = 22'b011_1011110101010100011;
                div_val= 22'b0000_010001000111010100;
            end
            10'd448:begin
                sqrt_val = 22'b011_1011111001100110000;
                div_val= 22'b0000_010001000110000110;
            end
            10'd449:begin
                sqrt_val = 22'b011_1011111101110111011;
                div_val= 22'b0000_010001000100111000;
            end
            10'd450:begin
                sqrt_val = 22'b011_1100000010001000100;
                div_val= 22'b0000_010001000011101010;
            end
            10'd451:begin
                sqrt_val = 22'b011_1100000110011001010;
                div_val= 22'b0000_010001000010011101;
            end
            10'd452:begin
                sqrt_val = 22'b011_1100001010101001110;
                div_val= 22'b0000_010001000001010000;
            end
            10'd453:begin
                sqrt_val = 22'b011_1100001110111001111;
                div_val= 22'b0000_010001000000000011;
            end
            10'd454:begin
                sqrt_val = 22'b011_1100010011001001110;
                div_val= 22'b0000_010000111110110110;
            end
            10'd455:begin
                sqrt_val = 22'b011_1100010111011001010;
                div_val= 22'b0000_010000111101101010;
            end
            10'd456:begin
                sqrt_val = 22'b011_1100011011101000101;
                div_val= 22'b0000_010000111100011110;
            end
            10'd457:begin
                sqrt_val = 22'b011_1100011111110111100;
                div_val= 22'b0000_010000111011010010;
            end
            10'd458:begin
                sqrt_val = 22'b011_1100100100000110010;
                div_val= 22'b0000_010000111010000110;
            end
            10'd459:begin
                sqrt_val = 22'b011_1100101000010100101;
                div_val= 22'b0000_010000111000111011;
            end
            10'd460:begin
                sqrt_val = 22'b011_1100101100100010101;
                div_val= 22'b0000_010000110111110000;
            end
            10'd461:begin
                sqrt_val = 22'b011_1100110000110000100;
                div_val= 22'b0000_010000110110100101;
            end
            10'd462:begin
                sqrt_val = 22'b011_1100110100111110000;
                div_val= 22'b0000_010000110101011010;
            end
            10'd463:begin
                sqrt_val = 22'b011_1100111001001011001;
                div_val= 22'b0000_010000110100010000;
            end
            10'd464:begin
                sqrt_val = 22'b011_1100111101011000001;
                div_val= 22'b0000_010000110011000101;
            end
            10'd465:begin
                sqrt_val = 22'b011_1101000001100100110;
                div_val= 22'b0000_010000110001111011;
            end
            10'd466:begin
                sqrt_val = 22'b011_1101000101110001000;
                div_val= 22'b0000_010000110000110010;
            end
            10'd467:begin
                sqrt_val = 22'b011_1101001001111101001;
                div_val= 22'b0000_010000101111101000;
            end
            10'd468:begin
                sqrt_val = 22'b011_1101001110001000111;
                div_val= 22'b0000_010000101110011111;
            end
            10'd469:begin
                sqrt_val = 22'b011_1101010010010100011;
                div_val= 22'b0000_010000101101010110;
            end
            10'd470:begin
                sqrt_val = 22'b011_1101010110011111100;
                div_val= 22'b0000_010000101100001101;
            end
            10'd471:begin
                sqrt_val = 22'b011_1101011010101010011;
                div_val= 22'b0000_010000101011000101;
            end
            10'd472:begin
                sqrt_val = 22'b011_1101011110110101000;
                div_val= 22'b0000_010000101001111100;
            end
            10'd473:begin
                sqrt_val = 22'b011_1101100010111111011;
                div_val= 22'b0000_010000101000110100;
            end
            10'd474:begin
                sqrt_val = 22'b011_1101100111001001100;
                div_val= 22'b0000_010000100111101100;
            end
            10'd475:begin
                sqrt_val = 22'b011_1101101011010011010;
                div_val= 22'b0000_010000100110100101;
            end
            10'd476:begin
                sqrt_val = 22'b011_1101101111011100110;
                div_val= 22'b0000_010000100101011101;
            end
            10'd477:begin
                sqrt_val = 22'b011_1101110011100110000;
                div_val= 22'b0000_010000100100010110;
            end
            10'd478:begin
                sqrt_val = 22'b011_1101110111101110111;
                div_val= 22'b0000_010000100011001111;
            end
            10'd479:begin
                sqrt_val = 22'b011_1101111011110111101;
                div_val= 22'b0000_010000100010001001;
            end
            10'd480:begin
                sqrt_val = 22'b011_1110000000000000000;
                div_val= 22'b0000_010000100001000010;
            end
            10'd481:begin
                sqrt_val = 22'b011_1110000100001000001;
                div_val= 22'b0000_010000011111111100;
            end
            10'd482:begin
                sqrt_val = 22'b011_1110001000010000000;
                div_val= 22'b0000_010000011110110110;
            end
            10'd483:begin
                sqrt_val = 22'b011_1110001100010111100;
                div_val= 22'b0000_010000011101110000;
            end
            10'd484:begin
                sqrt_val = 22'b011_1110010000011110111;
                div_val= 22'b0000_010000011100101010;
            end
            10'd485:begin
                sqrt_val = 22'b011_1110010100100101111;
                div_val= 22'b0000_010000011011100101;
            end
            10'd486:begin
                sqrt_val = 22'b011_1110011000101100101;
                div_val= 22'b0000_010000011010100000;
            end
            10'd487:begin
                sqrt_val = 22'b011_1110011100110011001;
                div_val= 22'b0000_010000011001011011;
            end
            10'd488:begin
                sqrt_val = 22'b011_1110100000111001011;
                div_val= 22'b0000_010000011000010110;
            end
            10'd489:begin
                sqrt_val = 22'b011_1110100100111111010;
                div_val= 22'b0000_010000010111010001;
            end
            10'd490:begin
                sqrt_val = 22'b011_1110101001000101000;
                div_val= 22'b0000_010000010110001101;
            end
            10'd491:begin
                sqrt_val = 22'b011_1110101101001010011;
                div_val= 22'b0000_010000010101001001;
            end
            10'd492:begin
                sqrt_val = 22'b011_1110110001001111100;
                div_val= 22'b0000_010000010100000101;
            end
            10'd493:begin
                sqrt_val = 22'b011_1110110101010100011;
                div_val= 22'b0000_010000010011000001;
            end
            10'd494:begin
                sqrt_val = 22'b011_1110111001011001000;
                div_val= 22'b0000_010000010001111110;
            end
            10'd495:begin
                sqrt_val = 22'b011_1110111101011101011;
                div_val= 22'b0000_010000010000111010;
            end
            10'd496:begin
                sqrt_val = 22'b011_1111000001100001100;
                div_val= 22'b0000_010000001111110111;
            end
            10'd497:begin
                sqrt_val = 22'b011_1111000101100101011;
                div_val= 22'b0000_010000001110110100;
            end
            10'd498:begin
                sqrt_val = 22'b011_1111001001101000111;
                div_val= 22'b0000_010000001101110001;
            end
            10'd499:begin
                sqrt_val = 22'b011_1111001101101100010;
                div_val= 22'b0000_010000001100101111;
            end
            10'd500:begin
                sqrt_val = 22'b011_1111010001101111010;
                div_val= 22'b0000_010000001011101101;
            end
            10'd501:begin
                sqrt_val = 22'b011_1111010101110010001;
                div_val= 22'b0000_010000001010101011;
            end
            10'd502:begin
                sqrt_val = 22'b011_1111011001110100101;
                div_val= 22'b0000_010000001001101001;
            end
            10'd503:begin
                sqrt_val = 22'b011_1111011101110110111;
                div_val= 22'b0000_010000001000100111;
            end
            10'd504:begin
                sqrt_val = 22'b011_1111100001111000111;
                div_val= 22'b0000_010000000111100101;
            end
            10'd505:begin
                sqrt_val = 22'b011_1111100101111010101;
                div_val= 22'b0000_010000000110100100;
            end
            10'd506:begin
                sqrt_val = 22'b011_1111101001111100010;
                div_val= 22'b0000_010000000101100011;
            end
            10'd507:begin
                sqrt_val = 22'b011_1111101101111101100;
                div_val= 22'b0000_010000000100100010;
            end
            10'd508:begin
                sqrt_val = 22'b011_1111110001111110100;
                div_val= 22'b0000_010000000011100001;
            end
            10'd509:begin
                sqrt_val = 22'b011_1111110101111111010;
                div_val= 22'b0000_010000000010100001;
            end
            10'd510:begin
                sqrt_val = 22'b011_1111111001111111110;
                div_val= 22'b0000_010000000001100000;
            end
            10'd511:begin
                sqrt_val = 22'b011_1111111110000000000;
                div_val= 22'b0000_010000000000100000;
            end
            10'd512:begin
                sqrt_val = 22'b100_0000000010000000000;
                div_val= 22'b0000_001111111111100000;
            end
            10'd513:begin
                sqrt_val = 22'b100_0000000101111111110;
                div_val= 22'b0000_001111111110100000;
            end
            10'd514:begin
                sqrt_val = 22'b100_0000001001111111010;
                div_val= 22'b0000_001111111101100001;
            end
            10'd515:begin
                sqrt_val = 22'b100_0000001101111110100;
                div_val= 22'b0000_001111111100100001;
            end
            10'd516:begin
                sqrt_val = 22'b100_0000010001111101100;
                div_val= 22'b0000_001111111011100010;
            end
            10'd517:begin
                sqrt_val = 22'b100_0000010101111100010;
                div_val= 22'b0000_001111111010100011;
            end
            10'd518:begin
                sqrt_val = 22'b100_0000011001111010110;
                div_val= 22'b0000_001111111001100100;
            end
            10'd519:begin
                sqrt_val = 22'b100_0000011101111001000;
                div_val= 22'b0000_001111111000100101;
            end
            10'd520:begin
                sqrt_val = 22'b100_0000100001110111000;
                div_val= 22'b0000_001111110111100111;
            end
            10'd521:begin
                sqrt_val = 22'b100_0000100101110100111;
                div_val= 22'b0000_001111110110101000;
            end
            10'd522:begin
                sqrt_val = 22'b100_0000101001110010011;
                div_val= 22'b0000_001111110101101010;
            end
            10'd523:begin
                sqrt_val = 22'b100_0000101101101111101;
                div_val= 22'b0000_001111110100101100;
            end
            10'd524:begin
                sqrt_val = 22'b100_0000110001101100110;
                div_val= 22'b0000_001111110011101110;
            end
            10'd525:begin
                sqrt_val = 22'b100_0000110101101001100;
                div_val= 22'b0000_001111110010110001;
            end
            10'd526:begin
                sqrt_val = 22'b100_0000111001100110001;
                div_val= 22'b0000_001111110001110011;
            end
            10'd527:begin
                sqrt_val = 22'b100_0000111101100010011;
                div_val= 22'b0000_001111110000110110;
            end
            10'd528:begin
                sqrt_val = 22'b100_0001000001011110100;
                div_val= 22'b0000_001111101111111001;
            end
            10'd529:begin
                sqrt_val = 22'b100_0001000101011010011;
                div_val= 22'b0000_001111101110111100;
            end
            10'd530:begin
                sqrt_val = 22'b100_0001001001010110000;
                div_val= 22'b0000_001111101101111111;
            end
            10'd531:begin
                sqrt_val = 22'b100_0001001101010001011;
                div_val= 22'b0000_001111101101000011;
            end
            10'd532:begin
                sqrt_val = 22'b100_0001010001001100100;
                div_val= 22'b0000_001111101100000110;
            end
            10'd533:begin
                sqrt_val = 22'b100_0001010101000111011;
                div_val= 22'b0000_001111101011001010;
            end
            10'd534:begin
                sqrt_val = 22'b100_0001011001000010001;
                div_val= 22'b0000_001111101010001110;
            end
            10'd535:begin
                sqrt_val = 22'b100_0001011100111100100;
                div_val= 22'b0000_001111101001010010;
            end
            10'd536:begin
                sqrt_val = 22'b100_0001100000110110110;
                div_val= 22'b0000_001111101000010110;
            end
            10'd537:begin
                sqrt_val = 22'b100_0001100100110000101;
                div_val= 22'b0000_001111100111011011;
            end
            10'd538:begin
                sqrt_val = 22'b100_0001101000101010011;
                div_val= 22'b0000_001111100110011111;
            end
            10'd539:begin
                sqrt_val = 22'b100_0001101100100011111;
                div_val= 22'b0000_001111100101100100;
            end
            10'd540:begin
                sqrt_val = 22'b100_0001110000011101010;
                div_val= 22'b0000_001111100100101001;
            end
            10'd541:begin
                sqrt_val = 22'b100_0001110100010110010;
                div_val= 22'b0000_001111100011101110;
            end
            10'd542:begin
                sqrt_val = 22'b100_0001111000001111000;
                div_val= 22'b0000_001111100010110011;
            end
            10'd543:begin
                sqrt_val = 22'b100_0001111100000111101;
                div_val= 22'b0000_001111100001111000;
            end
            10'd544:begin
                sqrt_val = 22'b100_0010000000000000000;
                div_val= 22'b0000_001111100000111110;
            end
            10'd545:begin
                sqrt_val = 22'b100_0010000011111000001;
                div_val= 22'b0000_001111100000000100;
            end
            10'd546:begin
                sqrt_val = 22'b100_0010000111110000000;
                div_val= 22'b0000_001111011111001010;
            end
            10'd547:begin
                sqrt_val = 22'b100_0010001011100111110;
                div_val= 22'b0000_001111011110010000;
            end
            10'd548:begin
                sqrt_val = 22'b100_0010001111011111001;
                div_val= 22'b0000_001111011101010110;
            end
            10'd549:begin
                sqrt_val = 22'b100_0010010011010110011;
                div_val= 22'b0000_001111011100011100;
            end
            10'd550:begin
                sqrt_val = 22'b100_0010010111001101011;
                div_val= 22'b0000_001111011011100011;
            end
            10'd551:begin
                sqrt_val = 22'b100_0010011011000100001;
                div_val= 22'b0000_001111011010101001;
            end
            10'd552:begin
                sqrt_val = 22'b100_0010011110111010110;
                div_val= 22'b0000_001111011001110000;
            end
            10'd553:begin
                sqrt_val = 22'b100_0010100010110001000;
                div_val= 22'b0000_001111011000110111;
            end
            10'd554:begin
                sqrt_val = 22'b100_0010100110100111001;
                div_val= 22'b0000_001111010111111110;
            end
            10'd555:begin
                sqrt_val = 22'b100_0010101010011101000;
                div_val= 22'b0000_001111010111000110;
            end
            10'd556:begin
                sqrt_val = 22'b100_0010101110010010101;
                div_val= 22'b0000_001111010110001101;
            end
            10'd557:begin
                sqrt_val = 22'b100_0010110010001000001;
                div_val= 22'b0000_001111010101010101;
            end
            10'd558:begin
                sqrt_val = 22'b100_0010110101111101011;
                div_val= 22'b0000_001111010100011100;
            end
            10'd559:begin
                sqrt_val = 22'b100_0010111001110010011;
                div_val= 22'b0000_001111010011100100;
            end
            10'd560:begin
                sqrt_val = 22'b100_0010111101100111001;
                div_val= 22'b0000_001111010010101100;
            end
            10'd561:begin
                sqrt_val = 22'b100_0011000001011011101;
                div_val= 22'b0000_001111010001110101;
            end
            10'd562:begin
                sqrt_val = 22'b100_0011000101010000000;
                div_val= 22'b0000_001111010000111101;
            end
            10'd563:begin
                sqrt_val = 22'b100_0011001001000100001;
                div_val= 22'b0000_001111010000000101;
            end
            10'd564:begin
                sqrt_val = 22'b100_0011001100111000001;
                div_val= 22'b0000_001111001111001110;
            end
            10'd565:begin
                sqrt_val = 22'b100_0011010000101011110;
                div_val= 22'b0000_001111001110010111;
            end
            10'd566:begin
                sqrt_val = 22'b100_0011010100011111010;
                div_val= 22'b0000_001111001101100000;
            end
            10'd567:begin
                sqrt_val = 22'b100_0011011000010010100;
                div_val= 22'b0000_001111001100101001;
            end
            10'd568:begin
                sqrt_val = 22'b100_0011011100000101101;
                div_val= 22'b0000_001111001011110010;
            end
            10'd569:begin
                sqrt_val = 22'b100_0011011111111000011;
                div_val= 22'b0000_001111001010111100;
            end
            10'd570:begin
                sqrt_val = 22'b100_0011100011101011000;
                div_val= 22'b0000_001111001010000101;
            end
            10'd571:begin
                sqrt_val = 22'b100_0011100111011101100;
                div_val= 22'b0000_001111001001001111;
            end
            10'd572:begin
                sqrt_val = 22'b100_0011101011001111101;
                div_val= 22'b0000_001111001000011001;
            end
            10'd573:begin
                sqrt_val = 22'b100_0011101111000001101;
                div_val= 22'b0000_001111000111100010;
            end
            10'd574:begin
                sqrt_val = 22'b100_0011110010110011011;
                div_val= 22'b0000_001111000110101101;
            end
            10'd575:begin
                sqrt_val = 22'b100_0011110110100101000;
                div_val= 22'b0000_001111000101110111;
            end
            10'd576:begin
                sqrt_val = 22'b100_0011111010010110011;
                div_val= 22'b0000_001111000101000001;
            end
            10'd577:begin
                sqrt_val = 22'b100_0011111110000111100;
                div_val= 22'b0000_001111000100001100;
            end
            10'd578:begin
                sqrt_val = 22'b100_0100000001111000100;
                div_val= 22'b0000_001111000011010110;
            end
            10'd579:begin
                sqrt_val = 22'b100_0100000101101001001;
                div_val= 22'b0000_001111000010100001;
            end
            10'd580:begin
                sqrt_val = 22'b100_0100001001011001110;
                div_val= 22'b0000_001111000001101100;
            end
            10'd581:begin
                sqrt_val = 22'b100_0100001101001010000;
                div_val= 22'b0000_001111000000110111;
            end
            10'd582:begin
                sqrt_val = 22'b100_0100010000111010001;
                div_val= 22'b0000_001111000000000010;
            end
            10'd583:begin
                sqrt_val = 22'b100_0100010100101010000;
                div_val= 22'b0000_001110111111001110;
            end
            10'd584:begin
                sqrt_val = 22'b100_0100011000011001110;
                div_val= 22'b0000_001110111110011001;
            end
            10'd585:begin
                sqrt_val = 22'b100_0100011100001001010;
                div_val= 22'b0000_001110111101100101;
            end
            10'd586:begin
                sqrt_val = 22'b100_0100011111111000100;
                div_val= 22'b0000_001110111100110000;
            end
            10'd587:begin
                sqrt_val = 22'b100_0100100011100111101;
                div_val= 22'b0000_001110111011111100;
            end
            10'd588:begin
                sqrt_val = 22'b100_0100100111010110100;
                div_val= 22'b0000_001110111011001000;
            end
            10'd589:begin
                sqrt_val = 22'b100_0100101011000101001;
                div_val= 22'b0000_001110111010010100;
            end
            10'd590:begin
                sqrt_val = 22'b100_0100101110110011101;
                div_val= 22'b0000_001110111001100001;
            end
            10'd591:begin
                sqrt_val = 22'b100_0100110010100001111;
                div_val= 22'b0000_001110111000101101;
            end
            10'd592:begin
                sqrt_val = 22'b100_0100110110010000000;
                div_val= 22'b0000_001110110111111010;
            end
            10'd593:begin
                sqrt_val = 22'b100_0100111001111101111;
                div_val= 22'b0000_001110110111000110;
            end
            10'd594:begin
                sqrt_val = 22'b100_0100111101101011100;
                div_val= 22'b0000_001110110110010011;
            end
            10'd595:begin
                sqrt_val = 22'b100_0101000001011001000;
                div_val= 22'b0000_001110110101100000;
            end
            10'd596:begin
                sqrt_val = 22'b100_0101000101000110010;
                div_val= 22'b0000_001110110100101101;
            end
            10'd597:begin
                sqrt_val = 22'b100_0101001000110011011;
                div_val= 22'b0000_001110110011111010;
            end
            10'd598:begin
                sqrt_val = 22'b100_0101001100100000010;
                div_val= 22'b0000_001110110011000111;
            end
            10'd599:begin
                sqrt_val = 22'b100_0101010000001101000;
                div_val= 22'b0000_001110110010010101;
            end
            10'd600:begin
                sqrt_val = 22'b100_0101010011111001011;
                div_val= 22'b0000_001110110001100010;
            end
            10'd601:begin
                sqrt_val = 22'b100_0101010111100101110;
                div_val= 22'b0000_001110110000110000;
            end
            10'd602:begin
                sqrt_val = 22'b100_0101011011010001110;
                div_val= 22'b0000_001110101111111110;
            end
            10'd603:begin
                sqrt_val = 22'b100_0101011110111101110;
                div_val= 22'b0000_001110101111001100;
            end
            10'd604:begin
                sqrt_val = 22'b100_0101100010101001011;
                div_val= 22'b0000_001110101110011010;
            end
            10'd605:begin
                sqrt_val = 22'b100_0101100110010100111;
                div_val= 22'b0000_001110101101101000;
            end
            10'd606:begin
                sqrt_val = 22'b100_0101101010000000010;
                div_val= 22'b0000_001110101100110110;
            end
            10'd607:begin
                sqrt_val = 22'b100_0101101101101011011;
                div_val= 22'b0000_001110101100000101;
            end
            10'd608:begin
                sqrt_val = 22'b100_0101110001010110010;
                div_val= 22'b0000_001110101011010011;
            end
            10'd609:begin
                sqrt_val = 22'b100_0101110101000001000;
                div_val= 22'b0000_001110101010100010;
            end
            10'd610:begin
                sqrt_val = 22'b100_0101111000101011100;
                div_val= 22'b0000_001110101001110001;
            end
            10'd611:begin
                sqrt_val = 22'b100_0101111100010101111;
                div_val= 22'b0000_001110101001000000;
            end
            10'd612:begin
                sqrt_val = 22'b100_0110000000000000000;
                div_val= 22'b0000_001110101000001111;
            end
            10'd613:begin
                sqrt_val = 22'b100_0110000011101010000;
                div_val= 22'b0000_001110100111011110;
            end
            10'd614:begin
                sqrt_val = 22'b100_0110000111010011110;
                div_val= 22'b0000_001110100110101101;
            end
            10'd615:begin
                sqrt_val = 22'b100_0110001010111101011;
                div_val= 22'b0000_001110100101111100;
            end
            10'd616:begin
                sqrt_val = 22'b100_0110001110100110110;
                div_val= 22'b0000_001110100101001100;
            end
            10'd617:begin
                sqrt_val = 22'b100_0110010010001111111;
                div_val= 22'b0000_001110100100011100;
            end
            10'd618:begin
                sqrt_val = 22'b100_0110010101111000111;
                div_val= 22'b0000_001110100011101011;
            end
            10'd619:begin
                sqrt_val = 22'b100_0110011001100001110;
                div_val= 22'b0000_001110100010111011;
            end
            10'd620:begin
                sqrt_val = 22'b100_0110011101001010011;
                div_val= 22'b0000_001110100010001011;
            end
            10'd621:begin
                sqrt_val = 22'b100_0110100000110010111;
                div_val= 22'b0000_001110100001011011;
            end
            10'd622:begin
                sqrt_val = 22'b100_0110100100011011001;
                div_val= 22'b0000_001110100000101011;
            end
            10'd623:begin
                sqrt_val = 22'b100_0110101000000011001;
                div_val= 22'b0000_001110011111111100;
            end
            10'd624:begin
                sqrt_val = 22'b100_0110101011101011000;
                div_val= 22'b0000_001110011111001100;
            end
            10'd625:begin
                sqrt_val = 22'b100_0110101111010010110;
                div_val= 22'b0000_001110011110011101;
            end
            10'd626:begin
                sqrt_val = 22'b100_0110110010111010010;
                div_val= 22'b0000_001110011101101101;
            end
            10'd627:begin
                sqrt_val = 22'b100_0110110110100001101;
                div_val= 22'b0000_001110011100111110;
            end
            10'd628:begin
                sqrt_val = 22'b100_0110111010001000110;
                div_val= 22'b0000_001110011100001111;
            end
            10'd629:begin
                sqrt_val = 22'b100_0110111101101111110;
                div_val= 22'b0000_001110011011100000;
            end
            10'd630:begin
                sqrt_val = 22'b100_0111000001010110100;
                div_val= 22'b0000_001110011010110001;
            end
            10'd631:begin
                sqrt_val = 22'b100_0111000100111101001;
                div_val= 22'b0000_001110011010000010;
            end
            10'd632:begin
                sqrt_val = 22'b100_0111001000100011100;
                div_val= 22'b0000_001110011001010100;
            end
            10'd633:begin
                sqrt_val = 22'b100_0111001100001001110;
                div_val= 22'b0000_001110011000100101;
            end
            10'd634:begin
                sqrt_val = 22'b100_0111001111101111111;
                div_val= 22'b0000_001110010111110111;
            end
            10'd635:begin
                sqrt_val = 22'b100_0111010011010101110;
                div_val= 22'b0000_001110010111001000;
            end
            10'd636:begin
                sqrt_val = 22'b100_0111010110111011011;
                div_val= 22'b0000_001110010110011010;
            end
            10'd637:begin
                sqrt_val = 22'b100_0111011010100000111;
                div_val= 22'b0000_001110010101101100;
            end
            10'd638:begin
                sqrt_val = 22'b100_0111011110000110010;
                div_val= 22'b0000_001110010100111110;
            end
            10'd639:begin
                sqrt_val = 22'b100_0111100001101011011;
                div_val= 22'b0000_001110010100010000;
            end
            10'd640:begin
                sqrt_val = 22'b100_0111100101010000011;
                div_val= 22'b0000_001110010011100010;
            end
            10'd641:begin
                sqrt_val = 22'b100_0111101000110101001;
                div_val= 22'b0000_001110010010110101;
            end
            10'd642:begin
                sqrt_val = 22'b100_0111101100011001110;
                div_val= 22'b0000_001110010010000111;
            end
            10'd643:begin
                sqrt_val = 22'b100_0111101111111110010;
                div_val= 22'b0000_001110010001011010;
            end
            10'd644:begin
                sqrt_val = 22'b100_0111110011100010100;
                div_val= 22'b0000_001110010000101100;
            end
            10'd645:begin
                sqrt_val = 22'b100_0111110111000110100;
                div_val= 22'b0000_001110001111111111;
            end
            10'd646:begin
                sqrt_val = 22'b100_0111111010101010100;
                div_val= 22'b0000_001110001111010010;
            end
            10'd647:begin
                sqrt_val = 22'b100_0111111110001110010;
                div_val= 22'b0000_001110001110100101;
            end
            10'd648:begin
                sqrt_val = 22'b100_1000000001110001110;
                div_val= 22'b0000_001110001101111000;
            end
            10'd649:begin
                sqrt_val = 22'b100_1000000101010101001;
                div_val= 22'b0000_001110001101001011;
            end
            10'd650:begin
                sqrt_val = 22'b100_1000001000111000011;
                div_val= 22'b0000_001110001100011110;
            end
            10'd651:begin
                sqrt_val = 22'b100_1000001100011011011;
                div_val= 22'b0000_001110001011110010;
            end
            10'd652:begin
                sqrt_val = 22'b100_1000001111111110010;
                div_val= 22'b0000_001110001011000101;
            end
            10'd653:begin
                sqrt_val = 22'b100_1000010011100000111;
                div_val= 22'b0000_001110001010011001;
            end
            10'd654:begin
                sqrt_val = 22'b100_1000010111000011011;
                div_val= 22'b0000_001110001001101100;
            end
            10'd655:begin
                sqrt_val = 22'b100_1000011010100101110;
                div_val= 22'b0000_001110001001000000;
            end
            10'd656:begin
                sqrt_val = 22'b100_1000011110000111111;
                div_val= 22'b0000_001110001000010100;
            end
            10'd657:begin
                sqrt_val = 22'b100_1000100001101001111;
                div_val= 22'b0000_001110000111101000;
            end
            10'd658:begin
                sqrt_val = 22'b100_1000100101001011110;
                div_val= 22'b0000_001110000110111100;
            end
            10'd659:begin
                sqrt_val = 22'b100_1000101000101101011;
                div_val= 22'b0000_001110000110010000;
            end
            10'd660:begin
                sqrt_val = 22'b100_1000101100001110111;
                div_val= 22'b0000_001110000101100100;
            end
            10'd661:begin
                sqrt_val = 22'b100_1000101111110000001;
                div_val= 22'b0000_001110000100111001;
            end
            10'd662:begin
                sqrt_val = 22'b100_1000110011010001010;
                div_val= 22'b0000_001110000100001101;
            end
            10'd663:begin
                sqrt_val = 22'b100_1000110110110010010;
                div_val= 22'b0000_001110000011100010;
            end
            10'd664:begin
                sqrt_val = 22'b100_1000111010010011001;
                div_val= 22'b0000_001110000010110110;
            end
            10'd665:begin
                sqrt_val = 22'b100_1000111101110011110;
                div_val= 22'b0000_001110000010001011;
            end
            10'd666:begin
                sqrt_val = 22'b100_1001000001010100001;
                div_val= 22'b0000_001110000001100000;
            end
            10'd667:begin
                sqrt_val = 22'b100_1001000100110100100;
                div_val= 22'b0000_001110000000110101;
            end
            10'd668:begin
                sqrt_val = 22'b100_1001001000010100101;
                div_val= 22'b0000_001110000000001010;
            end
            10'd669:begin
                sqrt_val = 22'b100_1001001011110100100;
                div_val= 22'b0000_001101111111011111;
            end
            10'd670:begin
                sqrt_val = 22'b100_1001001111010100010;
                div_val= 22'b0000_001101111110110100;
            end
            10'd671:begin
                sqrt_val = 22'b100_1001010010110011111;
                div_val= 22'b0000_001101111110001010;
            end
            10'd672:begin
                sqrt_val = 22'b100_1001010110010011011;
                div_val= 22'b0000_001101111101011111;
            end
            10'd673:begin
                sqrt_val = 22'b100_1001011001110010101;
                div_val= 22'b0000_001101111100110101;
            end
            10'd674:begin
                sqrt_val = 22'b100_1001011101010001110;
                div_val= 22'b0000_001101111100001010;
            end
            10'd675:begin
                sqrt_val = 22'b100_1001100000110000110;
                div_val= 22'b0000_001101111011100000;
            end
            10'd676:begin
                sqrt_val = 22'b100_1001100100001111100;
                div_val= 22'b0000_001101111010110110;
            end
            10'd677:begin
                sqrt_val = 22'b100_1001100111101110001;
                div_val= 22'b0000_001101111010001100;
            end
            10'd678:begin
                sqrt_val = 22'b100_1001101011001100101;
                div_val= 22'b0000_001101111001100010;
            end
            10'd679:begin
                sqrt_val = 22'b100_1001101110101011000;
                div_val= 22'b0000_001101111000111000;
            end
            10'd680:begin
                sqrt_val = 22'b100_1001110010001001001;
                div_val= 22'b0000_001101111000001110;
            end
            10'd681:begin
                sqrt_val = 22'b100_1001110101100111000;
                div_val= 22'b0000_001101110111100100;
            end
            10'd682:begin
                sqrt_val = 22'b100_1001111001000100111;
                div_val= 22'b0000_001101110110111011;
            end
            10'd683:begin
                sqrt_val = 22'b100_1001111100100010100;
                div_val= 22'b0000_001101110110010001;
            end
            10'd684:begin
                sqrt_val = 22'b100_1010000000000000000;
                div_val= 22'b0000_001101110101101000;
            end
            10'd685:begin
                sqrt_val = 22'b100_1010000011011101011;
                div_val= 22'b0000_001101110100111110;
            end
            10'd686:begin
                sqrt_val = 22'b100_1010000110111010100;
                div_val= 22'b0000_001101110100010101;
            end
            10'd687:begin
                sqrt_val = 22'b100_1010001010010111100;
                div_val= 22'b0000_001101110011101100;
            end
            10'd688:begin
                sqrt_val = 22'b100_1010001101110100011;
                div_val= 22'b0000_001101110011000011;
            end
            10'd689:begin
                sqrt_val = 22'b100_1010010001010001000;
                div_val= 22'b0000_001101110010011010;
            end
            10'd690:begin
                sqrt_val = 22'b100_1010010100101101100;
                div_val= 22'b0000_001101110001110001;
            end
            10'd691:begin
                sqrt_val = 22'b100_1010011000001001111;
                div_val= 22'b0000_001101110001001000;
            end
            10'd692:begin
                sqrt_val = 22'b100_1010011011100110001;
                div_val= 22'b0000_001101110000011111;
            end
            10'd693:begin
                sqrt_val = 22'b100_1010011111000010001;
                div_val= 22'b0000_001101101111110111;
            end
            10'd694:begin
                sqrt_val = 22'b100_1010100010011110000;
                div_val= 22'b0000_001101101111001110;
            end
            10'd695:begin
                sqrt_val = 22'b100_1010100101111001110;
                div_val= 22'b0000_001101101110100110;
            end
            10'd696:begin
                sqrt_val = 22'b100_1010101001010101011;
                div_val= 22'b0000_001101101101111101;
            end
            10'd697:begin
                sqrt_val = 22'b100_1010101100110000110;
                div_val= 22'b0000_001101101101010101;
            end
            10'd698:begin
                sqrt_val = 22'b100_1010110000001100000;
                div_val= 22'b0000_001101101100101101;
            end
            10'd699:begin
                sqrt_val = 22'b100_1010110011100111001;
                div_val= 22'b0000_001101101100000101;
            end
            10'd700:begin
                sqrt_val = 22'b100_1010110111000010000;
                div_val= 22'b0000_001101101011011101;
            end
            10'd701:begin
                sqrt_val = 22'b100_1010111010011100110;
                div_val= 22'b0000_001101101010110101;
            end
            10'd702:begin
                sqrt_val = 22'b100_1010111101110111011;
                div_val= 22'b0000_001101101010001101;
            end
            10'd703:begin
                sqrt_val = 22'b100_1011000001010001111;
                div_val= 22'b0000_001101101001100101;
            end
            10'd704:begin
                sqrt_val = 22'b100_1011000100101100010;
                div_val= 22'b0000_001101101000111101;
            end
            10'd705:begin
                sqrt_val = 22'b100_1011001000000110011;
                div_val= 22'b0000_001101101000010110;
            end
            10'd706:begin
                sqrt_val = 22'b100_1011001011100000011;
                div_val= 22'b0000_001101100111101110;
            end
            10'd707:begin
                sqrt_val = 22'b100_1011001110111010010;
                div_val= 22'b0000_001101100111000111;
            end
            10'd708:begin
                sqrt_val = 22'b100_1011010010010100000;
                div_val= 22'b0000_001101100110100000;
            end
            10'd709:begin
                sqrt_val = 22'b100_1011010101101101100;
                div_val= 22'b0000_001101100101111000;
            end
            10'd710:begin
                sqrt_val = 22'b100_1011011001000110111;
                div_val= 22'b0000_001101100101010001;
            end
            10'd711:begin
                sqrt_val = 22'b100_1011011100100000001;
                div_val= 22'b0000_001101100100101010;
            end
            10'd712:begin
                sqrt_val = 22'b100_1011011111111001010;
                div_val= 22'b0000_001101100100000011;
            end
            10'd713:begin
                sqrt_val = 22'b100_1011100011010010001;
                div_val= 22'b0000_001101100011011100;
            end
            10'd714:begin
                sqrt_val = 22'b100_1011100110101010111;
                div_val= 22'b0000_001101100010110101;
            end
            10'd715:begin
                sqrt_val = 22'b100_1011101010000011101;
                div_val= 22'b0000_001101100010001110;
            end
            10'd716:begin
                sqrt_val = 22'b100_1011101101011100000;
                div_val= 22'b0000_001101100001101000;
            end
            10'd717:begin
                sqrt_val = 22'b100_1011110000110100011;
                div_val= 22'b0000_001101100001000001;
            end
            10'd718:begin
                sqrt_val = 22'b100_1011110100001100100;
                div_val= 22'b0000_001101100000011010;
            end
            10'd719:begin
                sqrt_val = 22'b100_1011110111100100101;
                div_val= 22'b0000_001101011111110100;
            end
            10'd720:begin
                sqrt_val = 22'b100_1011111010111100100;
                div_val= 22'b0000_001101011111001110;
            end
            10'd721:begin
                sqrt_val = 22'b100_1011111110010100010;
                div_val= 22'b0000_001101011110100111;
            end
            10'd722:begin
                sqrt_val = 22'b100_1100000001101011110;
                div_val= 22'b0000_001101011110000001;
            end
            10'd723:begin
                sqrt_val = 22'b100_1100000101000011010;
                div_val= 22'b0000_001101011101011011;
            end
            10'd724:begin
                sqrt_val = 22'b100_1100001000011010100;
                div_val= 22'b0000_001101011100110101;
            end
            10'd725:begin
                sqrt_val = 22'b100_1100001011110001101;
                div_val= 22'b0000_001101011100001111;
            end
            10'd726:begin
                sqrt_val = 22'b100_1100001111001000101;
                div_val= 22'b0000_001101011011101001;
            end
            10'd727:begin
                sqrt_val = 22'b100_1100010010011111011;
                div_val= 22'b0000_001101011011000011;
            end
            10'd728:begin
                sqrt_val = 22'b100_1100010101110110001;
                div_val= 22'b0000_001101011010011101;
            end
            10'd729:begin
                sqrt_val = 22'b100_1100011001001100101;
                div_val= 22'b0000_001101011001111000;
            end
            10'd730:begin
                sqrt_val = 22'b100_1100011100100011000;
                div_val= 22'b0000_001101011001010010;
            end
            10'd731:begin
                sqrt_val = 22'b100_1100011111111001010;
                div_val= 22'b0000_001101011000101101;
            end
            10'd732:begin
                sqrt_val = 22'b100_1100100011001111011;
                div_val= 22'b0000_001101011000000111;
            end
            10'd733:begin
                sqrt_val = 22'b100_1100100110100101011;
                div_val= 22'b0000_001101010111100010;
            end
            10'd734:begin
                sqrt_val = 22'b100_1100101001111011001;
                div_val= 22'b0000_001101010110111101;
            end
            10'd735:begin
                sqrt_val = 22'b100_1100101101010000111;
                div_val= 22'b0000_001101010110010111;
            end
            10'd736:begin
                sqrt_val = 22'b100_1100110000100110011;
                div_val= 22'b0000_001101010101110010;
            end
            10'd737:begin
                sqrt_val = 22'b100_1100110011111011110;
                div_val= 22'b0000_001101010101001101;
            end
            10'd738:begin
                sqrt_val = 22'b100_1100110111010001000;
                div_val= 22'b0000_001101010100101000;
            end
            10'd739:begin
                sqrt_val = 22'b100_1100111010100110000;
                div_val= 22'b0000_001101010100000011;
            end
            10'd740:begin
                sqrt_val = 22'b100_1100111101111011000;
                div_val= 22'b0000_001101010011011110;
            end
            10'd741:begin
                sqrt_val = 22'b100_1101000001001111110;
                div_val= 22'b0000_001101010010111010;
            end
            10'd742:begin
                sqrt_val = 22'b100_1101000100100100011;
                div_val= 22'b0000_001101010010010101;
            end
            10'd743:begin
                sqrt_val = 22'b100_1101000111111001000;
                div_val= 22'b0000_001101010001110000;
            end
            10'd744:begin
                sqrt_val = 22'b100_1101001011001101011;
                div_val= 22'b0000_001101010001001100;
            end
            10'd745:begin
                sqrt_val = 22'b100_1101001110100001100;
                div_val= 22'b0000_001101010000100111;
            end
            10'd746:begin
                sqrt_val = 22'b100_1101010001110101101;
                div_val= 22'b0000_001101010000000011;
            end
            10'd747:begin
                sqrt_val = 22'b100_1101010101001001101;
                div_val= 22'b0000_001101001111011111;
            end
            10'd748:begin
                sqrt_val = 22'b100_1101011000011101011;
                div_val= 22'b0000_001101001110111010;
            end
            10'd749:begin
                sqrt_val = 22'b100_1101011011110001000;
                div_val= 22'b0000_001101001110010110;
            end
            10'd750:begin
                sqrt_val = 22'b100_1101011111000100100;
                div_val= 22'b0000_001101001101110010;
            end
            10'd751:begin
                sqrt_val = 22'b100_1101100010010111111;
                div_val= 22'b0000_001101001101001110;
            end
            10'd752:begin
                sqrt_val = 22'b100_1101100101101011001;
                div_val= 22'b0000_001101001100101010;
            end
            10'd753:begin
                sqrt_val = 22'b100_1101101000111110010;
                div_val= 22'b0000_001101001100000110;
            end
            10'd754:begin
                sqrt_val = 22'b100_1101101100010001010;
                div_val= 22'b0000_001101001011100011;
            end
            10'd755:begin
                sqrt_val = 22'b100_1101101111100100000;
                div_val= 22'b0000_001101001010111111;
            end
            10'd756:begin
                sqrt_val = 22'b100_1101110010110110101;
                div_val= 22'b0000_001101001010011011;
            end
            10'd757:begin
                sqrt_val = 22'b100_1101110110001001010;
                div_val= 22'b0000_001101001001111000;
            end
            10'd758:begin
                sqrt_val = 22'b100_1101111001011011101;
                div_val= 22'b0000_001101001001010100;
            end
            10'd759:begin
                sqrt_val = 22'b100_1101111100101101111;
                div_val= 22'b0000_001101001000110001;
            end
            10'd760:begin
                sqrt_val = 22'b100_1110000000000000000;
                div_val= 22'b0000_001101001000001101;
            end
            10'd761:begin
                sqrt_val = 22'b100_1110000011010010000;
                div_val= 22'b0000_001101000111101010;
            end
            10'd762:begin
                sqrt_val = 22'b100_1110000110100011111;
                div_val= 22'b0000_001101000111000111;
            end
            10'd763:begin
                sqrt_val = 22'b100_1110001001110101100;
                div_val= 22'b0000_001101000110100011;
            end
            10'd764:begin
                sqrt_val = 22'b100_1110001101000111001;
                div_val= 22'b0000_001101000110000000;
            end
            10'd765:begin
                sqrt_val = 22'b100_1110010000011000100;
                div_val= 22'b0000_001101000101011101;
            end
            10'd766:begin
                sqrt_val = 22'b100_1110010011101001111;
                div_val= 22'b0000_001101000100111010;
            end
            10'd767:begin
                sqrt_val = 22'b100_1110010110111011000;
                div_val= 22'b0000_001101000100010111;
            end
            10'd768:begin
                sqrt_val = 22'b100_1110011010001100000;
                div_val= 22'b0000_001101000011110101;
            end
            10'd769:begin
                sqrt_val = 22'b100_1110011101011100111;
                div_val= 22'b0000_001101000011010010;
            end
            10'd770:begin
                sqrt_val = 22'b100_1110100000101101101;
                div_val= 22'b0000_001101000010101111;
            end
            10'd771:begin
                sqrt_val = 22'b100_1110100011111110010;
                div_val= 22'b0000_001101000010001100;
            end
            10'd772:begin
                sqrt_val = 22'b100_1110100111001110110;
                div_val= 22'b0000_001101000001101010;
            end
            10'd773:begin
                sqrt_val = 22'b100_1110101010011111001;
                div_val= 22'b0000_001101000001000111;
            end
            10'd774:begin
                sqrt_val = 22'b100_1110101101101111010;
                div_val= 22'b0000_001101000000100101;
            end
            10'd775:begin
                sqrt_val = 22'b100_1110110000111111011;
                div_val= 22'b0000_001101000000000011;
            end
            10'd776:begin
                sqrt_val = 22'b100_1110110100001111011;
                div_val= 22'b0000_001100111111100000;
            end
            10'd777:begin
                sqrt_val = 22'b100_1110110111011111001;
                div_val= 22'b0000_001100111110111110;
            end
            10'd778:begin
                sqrt_val = 22'b100_1110111010101110110;
                div_val= 22'b0000_001100111110011100;
            end
            10'd779:begin
                sqrt_val = 22'b100_1110111101111110011;
                div_val= 22'b0000_001100111101111010;
            end
            10'd780:begin
                sqrt_val = 22'b100_1111000001001101110;
                div_val= 22'b0000_001100111101011000;
            end
            10'd781:begin
                sqrt_val = 22'b100_1111000100011101000;
                div_val= 22'b0000_001100111100110110;
            end
            10'd782:begin
                sqrt_val = 22'b100_1111000111101100001;
                div_val= 22'b0000_001100111100010100;
            end
            10'd783:begin
                sqrt_val = 22'b100_1111001010111011010;
                div_val= 22'b0000_001100111011110010;
            end
            10'd784:begin
                sqrt_val = 22'b100_1111001110001010001;
                div_val= 22'b0000_001100111011010000;
            end
            10'd785:begin
                sqrt_val = 22'b100_1111010001011000111;
                div_val= 22'b0000_001100111010101110;
            end
            10'd786:begin
                sqrt_val = 22'b100_1111010100100111011;
                div_val= 22'b0000_001100111010001101;
            end
            10'd787:begin
                sqrt_val = 22'b100_1111010111110101111;
                div_val= 22'b0000_001100111001101011;
            end
            10'd788:begin
                sqrt_val = 22'b100_1111011011000100010;
                div_val= 22'b0000_001100111001001010;
            end
            10'd789:begin
                sqrt_val = 22'b100_1111011110010010100;
                div_val= 22'b0000_001100111000101000;
            end
            10'd790:begin
                sqrt_val = 22'b100_1111100001100000101;
                div_val= 22'b0000_001100111000000111;
            end
            10'd791:begin
                sqrt_val = 22'b100_1111100100101110100;
                div_val= 22'b0000_001100110111100110;
            end
            10'd792:begin
                sqrt_val = 22'b100_1111100111111100011;
                div_val= 22'b0000_001100110111000100;
            end
            10'd793:begin
                sqrt_val = 22'b100_1111101011001010001;
                div_val= 22'b0000_001100110110100011;
            end
            10'd794:begin
                sqrt_val = 22'b100_1111101110010111101;
                div_val= 22'b0000_001100110110000010;
            end
            10'd795:begin
                sqrt_val = 22'b100_1111110001100101001;
                div_val= 22'b0000_001100110101100001;
            end
            10'd796:begin
                sqrt_val = 22'b100_1111110100110010011;
                div_val= 22'b0000_001100110101000000;
            end
            10'd797:begin
                sqrt_val = 22'b100_1111110111111111101;
                div_val= 22'b0000_001100110100011111;
            end
            10'd798:begin
                sqrt_val = 22'b100_1111111011001100101;
                div_val= 22'b0000_001100110011111110;
            end
            10'd799:begin
                sqrt_val = 22'b100_1111111110011001101;
                div_val= 22'b0000_001100110011011101;
            end
            10'd800:begin
                sqrt_val = 22'b101_0000000001100110011;
                div_val= 22'b0000_001100110010111100;
            end
            10'd801:begin
                sqrt_val = 22'b101_0000000100110011000;
                div_val= 22'b0000_001100110010011100;
            end
            10'd802:begin
                sqrt_val = 22'b101_0000000111111111101;
                div_val= 22'b0000_001100110001111011;
            end
            10'd803:begin
                sqrt_val = 22'b101_0000001011001100000;
                div_val= 22'b0000_001100110001011010;
            end
            10'd804:begin
                sqrt_val = 22'b101_0000001110011000010;
                div_val= 22'b0000_001100110000111010;
            end
            10'd805:begin
                sqrt_val = 22'b101_0000010001100100100;
                div_val= 22'b0000_001100110000011001;
            end
            10'd806:begin
                sqrt_val = 22'b101_0000010100110000100;
                div_val= 22'b0000_001100101111111001;
            end
            10'd807:begin
                sqrt_val = 22'b101_0000010111111100011;
                div_val= 22'b0000_001100101111011001;
            end
            10'd808:begin
                sqrt_val = 22'b101_0000011011001000010;
                div_val= 22'b0000_001100101110111000;
            end
            10'd809:begin
                sqrt_val = 22'b101_0000011110010011111;
                div_val= 22'b0000_001100101110011000;
            end
            10'd810:begin
                sqrt_val = 22'b101_0000100001011111011;
                div_val= 22'b0000_001100101101111000;
            end
            10'd811:begin
                sqrt_val = 22'b101_0000100100101010110;
                div_val= 22'b0000_001100101101011000;
            end
            10'd812:begin
                sqrt_val = 22'b101_0000100111110110001;
                div_val= 22'b0000_001100101100111000;
            end
            10'd813:begin
                sqrt_val = 22'b101_0000101011000001010;
                div_val= 22'b0000_001100101100011000;
            end
            10'd814:begin
                sqrt_val = 22'b101_0000101110001100010;
                div_val= 22'b0000_001100101011111000;
            end
            10'd815:begin
                sqrt_val = 22'b101_0000110001010111001;
                div_val= 22'b0000_001100101011011000;
            end
            10'd816:begin
                sqrt_val = 22'b101_0000110100100010000;
                div_val= 22'b0000_001100101010111000;
            end
            10'd817:begin
                sqrt_val = 22'b101_0000110111101100101;
                div_val= 22'b0000_001100101010011001;
            end
            10'd818:begin
                sqrt_val = 22'b101_0000111010110111001;
                div_val= 22'b0000_001100101001111001;
            end
            10'd819:begin
                sqrt_val = 22'b101_0000111110000001100;
                div_val= 22'b0000_001100101001011001;
            end
            10'd820:begin
                sqrt_val = 22'b101_0001000001001011111;
                div_val= 22'b0000_001100101000111010;
            end
            10'd821:begin
                sqrt_val = 22'b101_0001000100010110000;
                div_val= 22'b0000_001100101000011010;
            end
            10'd822:begin
                sqrt_val = 22'b101_0001000111100000000;
                div_val= 22'b0000_001100100111111011;
            end
            10'd823:begin
                sqrt_val = 22'b101_0001001010101010000;
                div_val= 22'b0000_001100100111011011;
            end
            10'd824:begin
                sqrt_val = 22'b101_0001001101110011110;
                div_val= 22'b0000_001100100110111100;
            end
            10'd825:begin
                sqrt_val = 22'b101_0001010000111101011;
                div_val= 22'b0000_001100100110011101;
            end
            10'd826:begin
                sqrt_val = 22'b101_0001010100000111000;
                div_val= 22'b0000_001100100101111101;
            end
            10'd827:begin
                sqrt_val = 22'b101_0001010111010000011;
                div_val= 22'b0000_001100100101011110;
            end
            10'd828:begin
                sqrt_val = 22'b101_0001011010011001110;
                div_val= 22'b0000_001100100100111111;
            end
            10'd829:begin
                sqrt_val = 22'b101_0001011101100010111;
                div_val= 22'b0000_001100100100100000;
            end
            10'd830:begin
                sqrt_val = 22'b101_0001100000101100000;
                div_val= 22'b0000_001100100100000001;
            end
            10'd831:begin
                sqrt_val = 22'b101_0001100011110100111;
                div_val= 22'b0000_001100100011100010;
            end
            10'd832:begin
                sqrt_val = 22'b101_0001100110111101110;
                div_val= 22'b0000_001100100011000011;
            end
            10'd833:begin
                sqrt_val = 22'b101_0001101010000110100;
                div_val= 22'b0000_001100100010100100;
            end
            10'd834:begin
                sqrt_val = 22'b101_0001101101001111000;
                div_val= 22'b0000_001100100010000110;
            end
            10'd835:begin
                sqrt_val = 22'b101_0001110000010111100;
                div_val= 22'b0000_001100100001100111;
            end
            10'd836:begin
                sqrt_val = 22'b101_0001110011011111111;
                div_val= 22'b0000_001100100001001000;
            end
            10'd837:begin
                sqrt_val = 22'b101_0001110110101000000;
                div_val= 22'b0000_001100100000101010;
            end
            10'd838:begin
                sqrt_val = 22'b101_0001111001110000001;
                div_val= 22'b0000_001100100000001011;
            end
            10'd839:begin
                sqrt_val = 22'b101_0001111100111000001;
                div_val= 22'b0000_001100011111101101;
            end
            10'd840:begin
                sqrt_val = 22'b101_0010000000000000000;
                div_val= 22'b0000_001100011111001110;
            end
            10'd841:begin
                sqrt_val = 22'b101_0010000011000111110;
                div_val= 22'b0000_001100011110110000;
            end
            10'd842:begin
                sqrt_val = 22'b101_0010000110001111011;
                div_val= 22'b0000_001100011110010001;
            end
            10'd843:begin
                sqrt_val = 22'b101_0010001001010110111;
                div_val= 22'b0000_001100011101110011;
            end
            10'd844:begin
                sqrt_val = 22'b101_0010001100011110010;
                div_val= 22'b0000_001100011101010101;
            end
            10'd845:begin
                sqrt_val = 22'b101_0010001111100101100;
                div_val= 22'b0000_001100011100110111;
            end
            10'd846:begin
                sqrt_val = 22'b101_0010010010101100110;
                div_val= 22'b0000_001100011100011000;
            end
            10'd847:begin
                sqrt_val = 22'b101_0010010101110011110;
                div_val= 22'b0000_001100011011111010;
            end
            10'd848:begin
                sqrt_val = 22'b101_0010011000111010101;
                div_val= 22'b0000_001100011011011100;
            end
            10'd849:begin
                sqrt_val = 22'b101_0010011100000001100;
                div_val= 22'b0000_001100011010111110;
            end
            10'd850:begin
                sqrt_val = 22'b101_0010011111001000001;
                div_val= 22'b0000_001100011010100000;
            end
            10'd851:begin
                sqrt_val = 22'b101_0010100010001110110;
                div_val= 22'b0000_001100011010000011;
            end
            10'd852:begin
                sqrt_val = 22'b101_0010100101010101001;
                div_val= 22'b0000_001100011001100101;
            end
            10'd853:begin
                sqrt_val = 22'b101_0010101000011011100;
                div_val= 22'b0000_001100011001000111;
            end
            10'd854:begin
                sqrt_val = 22'b101_0010101011100001110;
                div_val= 22'b0000_001100011000101001;
            end
            10'd855:begin
                sqrt_val = 22'b101_0010101110100111111;
                div_val= 22'b0000_001100011000001100;
            end
            10'd856:begin
                sqrt_val = 22'b101_0010110001101101110;
                div_val= 22'b0000_001100010111101110;
            end
            10'd857:begin
                sqrt_val = 22'b101_0010110100110011101;
                div_val= 22'b0000_001100010111010000;
            end
            10'd858:begin
                sqrt_val = 22'b101_0010110111111001011;
                div_val= 22'b0000_001100010110110011;
            end
            10'd859:begin
                sqrt_val = 22'b101_0010111010111111001;
                div_val= 22'b0000_001100010110010110;
            end
            10'd860:begin
                sqrt_val = 22'b101_0010111110000100101;
                div_val= 22'b0000_001100010101111000;
            end
            10'd861:begin
                sqrt_val = 22'b101_0011000001001010000;
                div_val= 22'b0000_001100010101011011;
            end
            10'd862:begin
                sqrt_val = 22'b101_0011000100001111011;
                div_val= 22'b0000_001100010100111101;
            end
            10'd863:begin
                sqrt_val = 22'b101_0011000111010100100;
                div_val= 22'b0000_001100010100100000;
            end
            10'd864:begin
                sqrt_val = 22'b101_0011001010011001101;
                div_val= 22'b0000_001100010100000011;
            end
            10'd865:begin
                sqrt_val = 22'b101_0011001101011110100;
                div_val= 22'b0000_001100010011100110;
            end
            10'd866:begin
                sqrt_val = 22'b101_0011010000100011011;
                div_val= 22'b0000_001100010011001001;
            end
            10'd867:begin
                sqrt_val = 22'b101_0011010011101000001;
                div_val= 22'b0000_001100010010101100;
            end
            10'd868:begin
                sqrt_val = 22'b101_0011010110101100110;
                div_val= 22'b0000_001100010010001111;
            end
            10'd869:begin
                sqrt_val = 22'b101_0011011001110001010;
                div_val= 22'b0000_001100010001110010;
            end
            10'd870:begin
                sqrt_val = 22'b101_0011011100110101101;
                div_val= 22'b0000_001100010001010101;
            end
            10'd871:begin
                sqrt_val = 22'b101_0011011111111001111;
                div_val= 22'b0000_001100010000111000;
            end
            10'd872:begin
                sqrt_val = 22'b101_0011100010111110000;
                div_val= 22'b0000_001100010000011011;
            end
            10'd873:begin
                sqrt_val = 22'b101_0011100110000010001;
                div_val= 22'b0000_001100001111111111;
            end
            10'd874:begin
                sqrt_val = 22'b101_0011101001000110000;
                div_val= 22'b0000_001100001111100010;
            end
            10'd875:begin
                sqrt_val = 22'b101_0011101100001001111;
                div_val= 22'b0000_001100001111000101;
            end
            10'd876:begin
                sqrt_val = 22'b101_0011101111001101100;
                div_val= 22'b0000_001100001110101001;
            end
            10'd877:begin
                sqrt_val = 22'b101_0011110010010001001;
                div_val= 22'b0000_001100001110001100;
            end
            10'd878:begin
                sqrt_val = 22'b101_0011110101010100101;
                div_val= 22'b0000_001100001101110000;
            end
            10'd879:begin
                sqrt_val = 22'b101_0011111000011000000;
                div_val= 22'b0000_001100001101010011;
            end
            10'd880:begin
                sqrt_val = 22'b101_0011111011011011010;
                div_val= 22'b0000_001100001100110111;
            end
            10'd881:begin
                sqrt_val = 22'b101_0011111110011110100;
                div_val= 22'b0000_001100001100011010;
            end
            10'd882:begin
                sqrt_val = 22'b101_0100000001100001100;
                div_val= 22'b0000_001100001011111110;
            end
            10'd883:begin
                sqrt_val = 22'b101_0100000100100100100;
                div_val= 22'b0000_001100001011100010;
            end
            10'd884:begin
                sqrt_val = 22'b101_0100000111100111010;
                div_val= 22'b0000_001100001011000110;
            end
            10'd885:begin
                sqrt_val = 22'b101_0100001010101010000;
                div_val= 22'b0000_001100001010101001;
            end
            10'd886:begin
                sqrt_val = 22'b101_0100001101101100101;
                div_val= 22'b0000_001100001010001101;
            end
            10'd887:begin
                sqrt_val = 22'b101_0100010000101111001;
                div_val= 22'b0000_001100001001110001;
            end
            10'd888:begin
                sqrt_val = 22'b101_0100010011110001100;
                div_val= 22'b0000_001100001001010101;
            end
            10'd889:begin
                sqrt_val = 22'b101_0100010110110011110;
                div_val= 22'b0000_001100001000111001;
            end
            10'd890:begin
                sqrt_val = 22'b101_0100011001110101111;
                div_val= 22'b0000_001100001000011101;
            end
            10'd891:begin
                sqrt_val = 22'b101_0100011100111000000;
                div_val= 22'b0000_001100001000000001;
            end
            10'd892:begin
                sqrt_val = 22'b101_0100011111111010000;
                div_val= 22'b0000_001100000111100110;
            end
            10'd893:begin
                sqrt_val = 22'b101_0100100010111011110;
                div_val= 22'b0000_001100000111001010;
            end
            10'd894:begin
                sqrt_val = 22'b101_0100100101111101100;
                div_val= 22'b0000_001100000110101110;
            end
            10'd895:begin
                sqrt_val = 22'b101_0100101000111111001;
                div_val= 22'b0000_001100000110010010;
            end
            10'd896:begin
                sqrt_val = 22'b101_0100101100000000101;
                div_val= 22'b0000_001100000101110111;
            end
            10'd897:begin
                sqrt_val = 22'b101_0100101111000010001;
                div_val= 22'b0000_001100000101011011;
            end
            10'd898:begin
                sqrt_val = 22'b101_0100110010000011011;
                div_val= 22'b0000_001100000101000000;
            end
            10'd899:begin
                sqrt_val = 22'b101_0100110101000100101;
                div_val= 22'b0000_001100000100100100;
            end
            10'd900:begin
                sqrt_val = 22'b101_0100111000000101101;
                div_val= 22'b0000_001100000100001001;
            end
            10'd901:begin
                sqrt_val = 22'b101_0100111011000110101;
                div_val= 22'b0000_001100000011101101;
            end
            10'd902:begin
                sqrt_val = 22'b101_0100111110000111100;
                div_val= 22'b0000_001100000011010010;
            end
            10'd903:begin
                sqrt_val = 22'b101_0101000001001000010;
                div_val= 22'b0000_001100000010110111;
            end
            10'd904:begin
                sqrt_val = 22'b101_0101000100001000111;
                div_val= 22'b0000_001100000010011011;
            end
            10'd905:begin
                sqrt_val = 22'b101_0101000111001001100;
                div_val= 22'b0000_001100000010000000;
            end
            10'd906:begin
                sqrt_val = 22'b101_0101001010001001111;
                div_val= 22'b0000_001100000001100101;
            end
            10'd907:begin
                sqrt_val = 22'b101_0101001101001010010;
                div_val= 22'b0000_001100000001001010;
            end
            10'd908:begin
                sqrt_val = 22'b101_0101010000001010100;
                div_val= 22'b0000_001100000000101111;
            end
            10'd909:begin
                sqrt_val = 22'b101_0101010011001010101;
                div_val= 22'b0000_001100000000010100;
            end
            10'd910:begin
                sqrt_val = 22'b101_0101010110001010101;
                div_val= 22'b0000_001011111111111001;
            end
            10'd911:begin
                sqrt_val = 22'b101_0101011001001010101;
                div_val= 22'b0000_001011111111011110;
            end
            10'd912:begin
                sqrt_val = 22'b101_0101011100001010011;
                div_val= 22'b0000_001011111111000011;
            end
            10'd913:begin
                sqrt_val = 22'b101_0101011111001010001;
                div_val= 22'b0000_001011111110101000;
            end
            10'd914:begin
                sqrt_val = 22'b101_0101100010001001110;
                div_val= 22'b0000_001011111110001101;
            end
            10'd915:begin
                sqrt_val = 22'b101_0101100101001001010;
                div_val= 22'b0000_001011111101110010;
            end
            10'd916:begin
                sqrt_val = 22'b101_0101101000001000101;
                div_val= 22'b0000_001011111101010111;
            end
            10'd917:begin
                sqrt_val = 22'b101_0101101011000111111;
                div_val= 22'b0000_001011111100111101;
            end
            10'd918:begin
                sqrt_val = 22'b101_0101101110000111001;
                div_val= 22'b0000_001011111100100010;
            end
            10'd919:begin
                sqrt_val = 22'b101_0101110001000110001;
                div_val= 22'b0000_001011111100000111;
            end
            10'd920:begin
                sqrt_val = 22'b101_0101110100000101001;
                div_val= 22'b0000_001011111011101101;
            end
            10'd921:begin
                sqrt_val = 22'b101_0101110111000100000;
                div_val= 22'b0000_001011111011010010;
            end
            10'd922:begin
                sqrt_val = 22'b101_0101111010000010110;
                div_val= 22'b0000_001011111010111000;
            end
            10'd923:begin
                sqrt_val = 22'b101_0101111101000001011;
                div_val= 22'b0000_001011111010011101;
            end
            10'd924:begin
                sqrt_val = 22'b101_0110000000000000000;
                div_val= 22'b0000_001011111010000011;
            end
            10'd925:begin
                sqrt_val = 22'b101_0110000010111110100;
                div_val= 22'b0000_001011111001101001;
            end
            10'd926:begin
                sqrt_val = 22'b101_0110000101111100111;
                div_val= 22'b0000_001011111001001110;
            end
            10'd927:begin
                sqrt_val = 22'b101_0110001000111011001;
                div_val= 22'b0000_001011111000110100;
            end
            10'd928:begin
                sqrt_val = 22'b101_0110001011111001010;
                div_val= 22'b0000_001011111000011010;
            end
            10'd929:begin
                sqrt_val = 22'b101_0110001110110111010;
                div_val= 22'b0000_001011111000000000;
            end
            10'd930:begin
                sqrt_val = 22'b101_0110010001110101010;
                div_val= 22'b0000_001011110111100101;
            end
            10'd931:begin
                sqrt_val = 22'b101_0110010100110011001;
                div_val= 22'b0000_001011110111001011;
            end
            10'd932:begin
                sqrt_val = 22'b101_0110010111110000110;
                div_val= 22'b0000_001011110110110001;
            end
            10'd933:begin
                sqrt_val = 22'b101_0110011010101110100;
                div_val= 22'b0000_001011110110010111;
            end
            10'd934:begin
                sqrt_val = 22'b101_0110011101101100000;
                div_val= 22'b0000_001011110101111101;
            end
            10'd935:begin
                sqrt_val = 22'b101_0110100000101001011;
                div_val= 22'b0000_001011110101100011;
            end
            10'd936:begin
                sqrt_val = 22'b101_0110100011100110110;
                div_val= 22'b0000_001011110101001010;
            end
            10'd937:begin
                sqrt_val = 22'b101_0110100110100100000;
                div_val= 22'b0000_001011110100110000;
            end
            10'd938:begin
                sqrt_val = 22'b101_0110101001100001001;
                div_val= 22'b0000_001011110100010110;
            end
            10'd939:begin
                sqrt_val = 22'b101_0110101100011110001;
                div_val= 22'b0000_001011110011111100;
            end
            10'd940:begin
                sqrt_val = 22'b101_0110101111011011001;
                div_val= 22'b0000_001011110011100010;
            end
            10'd941:begin
                sqrt_val = 22'b101_0110110010011000000;
                div_val= 22'b0000_001011110011001001;
            end
            10'd942:begin
                sqrt_val = 22'b101_0110110101010100101;
                div_val= 22'b0000_001011110010101111;
            end
            10'd943:begin
                sqrt_val = 22'b101_0110111000010001010;
                div_val= 22'b0000_001011110010010101;
            end
            10'd944:begin
                sqrt_val = 22'b101_0110111011001101111;
                div_val= 22'b0000_001011110001111100;
            end
            10'd945:begin
                sqrt_val = 22'b101_0110111110001010010;
                div_val= 22'b0000_001011110001100010;
            end
            10'd946:begin
                sqrt_val = 22'b101_0111000001000110101;
                div_val= 22'b0000_001011110001001001;
            end
            10'd947:begin
                sqrt_val = 22'b101_0111000100000010111;
                div_val= 22'b0000_001011110000101111;
            end
            10'd948:begin
                sqrt_val = 22'b101_0111000110111111000;
                div_val= 22'b0000_001011110000010110;
            end
            10'd949:begin
                sqrt_val = 22'b101_0111001001111011000;
                div_val= 22'b0000_001011101111111101;
            end
            10'd950:begin
                sqrt_val = 22'b101_0111001100110111000;
                div_val= 22'b0000_001011101111100011;
            end
            10'd951:begin
                sqrt_val = 22'b101_0111001111110010110;
                div_val= 22'b0000_001011101111001010;
            end
            10'd952:begin
                sqrt_val = 22'b101_0111010010101110100;
                div_val= 22'b0000_001011101110110001;
            end
            10'd953:begin
                sqrt_val = 22'b101_0111010101101010001;
                div_val= 22'b0000_001011101110011000;
            end
            10'd954:begin
                sqrt_val = 22'b101_0111011000100101110;
                div_val= 22'b0000_001011101101111110;
            end
            10'd955:begin
                sqrt_val = 22'b101_0111011011100001001;
                div_val= 22'b0000_001011101101100101;
            end
            10'd956:begin
                sqrt_val = 22'b101_0111011110011100100;
                div_val= 22'b0000_001011101101001100;
            end
            10'd957:begin
                sqrt_val = 22'b101_0111100001010111110;
                div_val= 22'b0000_001011101100110011;
            end
            10'd958:begin
                sqrt_val = 22'b101_0111100100010010111;
                div_val= 22'b0000_001011101100011010;
            end
            10'd959:begin
                sqrt_val = 22'b101_0111100111001110000;
                div_val= 22'b0000_001011101100000001;
            end
            10'd960:begin
                sqrt_val = 22'b101_0111101010001000111;
                div_val= 22'b0000_001011101011101000;
            end
            10'd961:begin
                sqrt_val = 22'b101_0111101101000011110;
                div_val= 22'b0000_001011101011001111;
            end
            10'd962:begin
                sqrt_val = 22'b101_0111101111111110100;
                div_val= 22'b0000_001011101010110111;
            end
            10'd963:begin
                sqrt_val = 22'b101_0111110010111001010;
                div_val= 22'b0000_001011101010011110;
            end
            10'd964:begin
                sqrt_val = 22'b101_0111110101110011110;
                div_val= 22'b0000_001011101010000101;
            end
            10'd965:begin
                sqrt_val = 22'b101_0111111000101110010;
                div_val= 22'b0000_001011101001101100;
            end
            10'd966:begin
                sqrt_val = 22'b101_0111111011101000101;
                div_val= 22'b0000_001011101001010100;
            end
            10'd967:begin
                sqrt_val = 22'b101_0111111110100010111;
                div_val= 22'b0000_001011101000111011;
            end
            10'd968:begin
                sqrt_val = 22'b101_1000000001011101001;
                div_val= 22'b0000_001011101000100010;
            end
            10'd969:begin
                sqrt_val = 22'b101_1000000100010111001;
                div_val= 22'b0000_001011101000001010;
            end
            10'd970:begin
                sqrt_val = 22'b101_1000000111010001001;
                div_val= 22'b0000_001011100111110001;
            end
            10'd971:begin
                sqrt_val = 22'b101_1000001010001011000;
                div_val= 22'b0000_001011100111011001;
            end
            10'd972:begin
                sqrt_val = 22'b101_1000001101000100111;
                div_val= 22'b0000_001011100111000000;
            end
            10'd973:begin
                sqrt_val = 22'b101_1000001111111110100;
                div_val= 22'b0000_001011100110101000;
            end
            10'd974:begin
                sqrt_val = 22'b101_1000010010111000001;
                div_val= 22'b0000_001011100110001111;
            end
            10'd975:begin
                sqrt_val = 22'b101_1000010101110001101;
                div_val= 22'b0000_001011100101110111;
            end
            10'd976:begin
                sqrt_val = 22'b101_1000011000101011001;
                div_val= 22'b0000_001011100101011111;
            end
            10'd977:begin
                sqrt_val = 22'b101_1000011011100100011;
                div_val= 22'b0000_001011100101000110;
            end
            10'd978:begin
                sqrt_val = 22'b101_1000011110011101101;
                div_val= 22'b0000_001011100100101110;
            end
            10'd979:begin
                sqrt_val = 22'b101_1000100001010110110;
                div_val= 22'b0000_001011100100010110;
            end
            10'd980:begin
                sqrt_val = 22'b101_1000100100001111110;
                div_val= 22'b0000_001011100011111110;
            end
            10'd981:begin
                sqrt_val = 22'b101_1000100111001000110;
                div_val= 22'b0000_001011100011100110;
            end
            10'd982:begin
                sqrt_val = 22'b101_1000101010000001101;
                div_val= 22'b0000_001011100011001110;
            end
            10'd983:begin
                sqrt_val = 22'b101_1000101100111010011;
                div_val= 22'b0000_001011100010110101;
            end
            10'd984:begin
                sqrt_val = 22'b101_1000101111110011000;
                div_val= 22'b0000_001011100010011101;
            end
            10'd985:begin
                sqrt_val = 22'b101_1000110010101011101;
                div_val= 22'b0000_001011100010000101;
            end
            10'd986:begin
                sqrt_val = 22'b101_1000110101100100000;
                div_val= 22'b0000_001011100001101110;
            end
            10'd987:begin
                sqrt_val = 22'b101_1000111000011100100;
                div_val= 22'b0000_001011100001010110;
            end
            10'd988:begin
                sqrt_val = 22'b101_1000111011010100110;
                div_val= 22'b0000_001011100000111110;
            end
            10'd989:begin
                sqrt_val = 22'b101_1000111110001100111;
                div_val= 22'b0000_001011100000100110;
            end
            10'd990:begin
                sqrt_val = 22'b101_1001000001000101000;
                div_val= 22'b0000_001011100000001110;
            end
            10'd991:begin
                sqrt_val = 22'b101_1001000011111101000;
                div_val= 22'b0000_001011011111110110;
            end
            10'd992:begin
                sqrt_val = 22'b101_1001000110110101000;
                div_val= 22'b0000_001011011111011111;
            end
            10'd993:begin
                sqrt_val = 22'b101_1001001001101100110;
                div_val= 22'b0000_001011011111000111;
            end
            10'd994:begin
                sqrt_val = 22'b101_1001001100100100100;
                div_val= 22'b0000_001011011110101111;
            end
            10'd995:begin
                sqrt_val = 22'b101_1001001111011100001;
                div_val= 22'b0000_001011011110011000;
            end
            10'd996:begin
                sqrt_val = 22'b101_1001010010010011110;
                div_val= 22'b0000_001011011110000000;
            end
            10'd997:begin
                sqrt_val = 22'b101_1001010101001011001;
                div_val= 22'b0000_001011011101101000;
            end
            10'd998:begin
                sqrt_val = 22'b101_1001011000000010100;
                div_val= 22'b0000_001011011101010001;
            end
            10'd999:begin
                sqrt_val = 22'b101_1001011010111001110;
                div_val= 22'b0000_001011011100111001;
            end
            10'd1000:begin
                sqrt_val = 22'b101_1001011101110001000;
                div_val= 22'b0000_001011011100100010;
            end
            10'd1001:begin
                sqrt_val = 22'b101_1001100000101000000;
                div_val= 22'b0000_001011011100001011;
            end
            10'd1002:begin
                sqrt_val = 22'b101_1001100011011111000;
                div_val= 22'b0000_001011011011110011;
            end
            10'd1003:begin
                sqrt_val = 22'b101_1001100110010110000;
                div_val= 22'b0000_001011011011011100;
            end
            10'd1004:begin
                sqrt_val = 22'b101_1001101001001100110;
                div_val= 22'b0000_001011011011000101;
            end
            10'd1005:begin
                sqrt_val = 22'b101_1001101100000011100;
                div_val= 22'b0000_001011011010101101;
            end
            10'd1006:begin
                sqrt_val = 22'b101_1001101110111010001;
                div_val= 22'b0000_001011011010010110;
            end
            10'd1007:begin
                sqrt_val = 22'b101_1001110001110000101;
                div_val= 22'b0000_001011011001111111;
            end
            10'd1008:begin
                sqrt_val = 22'b101_1001110100100111001;
                div_val= 22'b0000_001011011001101000;
            end
            10'd1009:begin
                sqrt_val = 22'b101_1001110111011101100;
                div_val= 22'b0000_001011011001010001;
            end
            10'd1010:begin
                sqrt_val = 22'b101_1001111010010011110;
                div_val= 22'b0000_001011011000111001;
            end
            10'd1011:begin
                sqrt_val = 22'b101_1001111101001001111;
                div_val= 22'b0000_001011011000100010;
            end
            10'd1012:begin
                sqrt_val = 22'b101_1010000000000000000;
                div_val= 22'b0000_001011011000001011;
            end
            10'd1013:begin
                sqrt_val = 22'b101_1010000010110110000;
                div_val= 22'b0000_001011010111110100;
            end
            10'd1014:begin
                sqrt_val = 22'b101_1010000101101011111;
                div_val= 22'b0000_001011010111011101;
            end
            10'd1015:begin
                sqrt_val = 22'b101_1010001000100001110;
                div_val= 22'b0000_001011010111000110;
            end
            10'd1016:begin
                sqrt_val = 22'b101_1010001011010111100;
                div_val= 22'b0000_001011010110110000;
            end
            10'd1017:begin
                sqrt_val = 22'b101_1010001110001101001;
                div_val= 22'b0000_001011010110011001;
            end
            10'd1018:begin
                sqrt_val = 22'b101_1010010001000010101;
                div_val= 22'b0000_001011010110000010;
            end
            10'd1019:begin
                sqrt_val = 22'b101_1010010011111000001;
                div_val= 22'b0000_001011010101101011;
            end
            10'd1020:begin
                sqrt_val = 22'b101_1010010110101101100;
                div_val= 22'b0000_001011010101010100;
            end
            10'd1021:begin
                sqrt_val = 22'b101_1010011001100010110;
                div_val= 22'b0000_001011010100111110;
            end
            10'd1022:begin
                sqrt_val = 22'b101_1010011100011000000;
                div_val= 22'b0000_001011010100100111;
            end
            10'd1023:begin
                sqrt_val = 22'b101_1010011111001101001;
                div_val= 22'b0000_001011010100010000;
            end
            default:begin
                sqrt_val = 22'd0;
                div_val= 22'd0;
            end
        endcase
    end

endmodule

module complex_mul_48_40 ( 
    // input clk,
    // input rst,
    input [47:0] complex_in1,
    input [39:0] complex_in2,
    output [39:0] output_data//{{s,3,16},{s,3,16}}
);

    wire signed [20:0] tmp1,tmp2,tmp3,tmp4;
    wire signed [21:0] sum_real,sum_imag ;

    assign tmp1 =  $signed(complex_in1[23:13])*$signed(complex_in2[19:9]);//{s,1+3,11+9}
    assign tmp2 =  $signed(complex_in1[47:37])*$signed(complex_in2[39:29]);
    assign sum_real = $signed({tmp1[20],tmp1})-$signed({tmp2[20],tmp2});//{s,1+3+1,10+8}
    assign output_data[19:0] = {sum_real[20],sum_real[18:0]};

    assign tmp3 =  $signed(complex_in1[23:13])*$signed(complex_in2[39:29]);
    assign tmp4 =  $signed(complex_in1[47:37])*$signed(complex_in2[19:9]);
    assign sum_imag = $signed({tmp3[20],tmp3})+$signed({tmp4[20],tmp4}); //overflow?
    assign output_data[39:20] = {sum_imag[20],sum_imag[18:0]};

endmodule 

module complex_mul_40_40 ( 
    // input clk,
    // input rst,
    input [39:0] complex_in1,
    input [39:0] complex_in2,
    output [31:0] output_data//{{s,1,22},{s,1,22}}
);

    wire signed [18:0] tmp1,tmp2,tmp3,tmp4;
    wire signed [19:0] sum_real,sum_imag ;

    assign tmp1 =  $signed(complex_in1[19:10])*$signed(complex_in2[19:10]);   //{s1,8}{s3,6}={s4,14}
    assign tmp2 =  $signed(complex_in1[39:30])*$signed(complex_in2[39:30]);//{s,6,16}
    assign sum_real = $signed({tmp1[18],tmp1})-$signed({tmp2[18],tmp2});////{s,6+1,16} - {s,6+1,16}       {s5,14}
    assign output_data[15:0] = {sum_real[19],sum_real[14:0]};//{s,3,12}

    assign tmp3 =  $signed(complex_in1[19:10])*$signed(complex_in2[39:30]);
    assign tmp4 =  $signed(complex_in1[39:30])*$signed(complex_in2[19:10]);
    assign sum_imag = $signed({tmp3[18],tmp3})+$signed({tmp4[18],tmp4});//overflow?
    assign output_data[31:16] = {sum_imag[19],sum_imag[14:0]};



endmodule 
